/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Apr 23 17:02:10 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1347508157 */

module adder(A, B, is_subtract, result, carry, overflow_flag, negative);
   input [15:0]A;
   input [15:0]B;
   input is_subtract;
   output [15:0]result;
   output carry;
   output overflow_flag;
   output negative;

   wire n_0_0_0;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_54;
   wire n_0_0_51;
   wire n_0_0_50;
   wire n_0_0_48;
   wire n_0_0_46;
   wire n_0_0_44;
   wire n_0_0_43;
   wire n_0_0_41;
   wire n_0_0_39;
   wire n_0_0_37;
   wire n_0_0_36;
   wire n_0_0_34;
   wire n_0_0_32;
   wire n_0_0_30;
   wire n_0_0_29;
   wire n_0_0_27;
   wire n_0_0_25;
   wire n_0_0_23;
   wire n_0_0_22;
   wire n_0_0_20;
   wire n_0_0_18;
   wire n_0_0_16;
   wire n_0_0_15;
   wire n_0_0_13;
   wire n_0_0_11;
   wire n_0_0_9;
   wire n_0_0_3;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_6;
   wire n_0_0_8;
   wire n_0_0_10;
   wire n_0_0_12;
   wire n_0_0_14;
   wire n_0_0_17;
   wire n_0_0_19;
   wire n_0_0_21;
   wire n_0_0_24;
   wire n_0_0_26;
   wire n_0_0_28;
   wire n_0_0_31;
   wire n_0_0_33;
   wire n_0_0_35;
   wire n_0_0_38;
   wire n_0_0_40;
   wire n_0_0_42;
   wire n_0_0_45;
   wire n_0_0_47;
   wire n_0_0_49;
   wire n_0_0_52;
   wire n_0_0_7;
   wire n_0_0_53;
   wire n_0_0_55;
   wire n_0_0_5;
   wire n_0_0_4;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;

   XOR2_X1 i_0_0_0 (.A(B[15]), .B(is_subtract), .Z(n_0_0_0));
   XNOR2_X1 i_0_0_1 (.A(is_subtract), .B(A[0]), .ZN(n_0_0_60));
   OAI21_X1 i_0_0_2 (.A(n_0_0_5), .B1(n_0_0_4), .B2(is_subtract), .ZN(n_0_0_61));
   XNOR2_X1 i_0_0_3 (.A(n_0_0_60), .B(n_0_0_61), .ZN(result[0]));
   XNOR2_X1 i_0_0_4 (.A(n_0_0_3), .B(n_0_0_7), .ZN(result[1]));
   XOR2_X1 i_0_0_5 (.A(n_0_0_9), .B(n_0_0_11), .Z(result[2]));
   XOR2_X1 i_0_0_6 (.A(n_0_0_13), .B(n_0_0_15), .Z(result[3]));
   XOR2_X1 i_0_0_7 (.A(n_0_0_16), .B(n_0_0_18), .Z(result[4]));
   XOR2_X1 i_0_0_8 (.A(n_0_0_20), .B(n_0_0_22), .Z(result[5]));
   XOR2_X1 i_0_0_9 (.A(n_0_0_23), .B(n_0_0_25), .Z(result[6]));
   XOR2_X1 i_0_0_10 (.A(n_0_0_27), .B(n_0_0_29), .Z(result[7]));
   XOR2_X1 i_0_0_11 (.A(n_0_0_30), .B(n_0_0_32), .Z(result[8]));
   XOR2_X1 i_0_0_12 (.A(n_0_0_34), .B(n_0_0_36), .Z(result[9]));
   XOR2_X1 i_0_0_13 (.A(n_0_0_39), .B(n_0_0_37), .Z(result[10]));
   XOR2_X1 i_0_0_14 (.A(n_0_0_41), .B(n_0_0_43), .Z(result[11]));
   XOR2_X1 i_0_0_15 (.A(n_0_0_46), .B(n_0_0_44), .Z(result[12]));
   XOR2_X1 i_0_0_16 (.A(n_0_0_48), .B(n_0_0_50), .Z(result[13]));
   XNOR2_X1 i_0_0_17 (.A(n_0_0_51), .B(n_0_0_54), .ZN(result[14]));
   NOR2_X1 i_0_0_18 (.A1(n_0_0_127), .A2(n_0_0_130), .ZN(n_0_0_54));
   NAND2_X1 i_0_0_19 (.A1(n_0_0_24), .A2(n_0_0_124), .ZN(n_0_0_51));
   AND2_X1 i_0_0_20 (.A1(n_0_0_124), .A2(n_0_0_123), .ZN(n_0_0_50));
   NOR2_X1 i_0_0_21 (.A1(n_0_0_26), .A2(n_0_0_117), .ZN(n_0_0_48));
   OR2_X1 i_0_0_22 (.A1(n_0_0_117), .A2(n_0_0_116), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_23 (.A1(n_0_0_28), .A2(n_0_0_113), .ZN(n_0_0_44));
   AND2_X1 i_0_0_24 (.A1(n_0_0_113), .A2(n_0_0_112), .ZN(n_0_0_43));
   NOR2_X1 i_0_0_25 (.A1(n_0_0_31), .A2(n_0_0_107), .ZN(n_0_0_41));
   OR2_X1 i_0_0_26 (.A1(n_0_0_107), .A2(n_0_0_106), .ZN(n_0_0_39));
   NAND2_X1 i_0_0_27 (.A1(n_0_0_33), .A2(n_0_0_103), .ZN(n_0_0_37));
   AND2_X1 i_0_0_28 (.A1(n_0_0_103), .A2(n_0_0_102), .ZN(n_0_0_36));
   NOR2_X1 i_0_0_29 (.A1(n_0_0_35), .A2(n_0_0_97), .ZN(n_0_0_34));
   OR2_X1 i_0_0_30 (.A1(n_0_0_97), .A2(n_0_0_96), .ZN(n_0_0_32));
   NAND2_X1 i_0_0_31 (.A1(n_0_0_38), .A2(n_0_0_93), .ZN(n_0_0_30));
   AND2_X1 i_0_0_32 (.A1(n_0_0_93), .A2(n_0_0_92), .ZN(n_0_0_29));
   NOR2_X1 i_0_0_33 (.A1(n_0_0_40), .A2(n_0_0_87), .ZN(n_0_0_27));
   OR2_X1 i_0_0_34 (.A1(n_0_0_87), .A2(n_0_0_86), .ZN(n_0_0_25));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_42), .A2(n_0_0_83), .ZN(n_0_0_23));
   AND2_X1 i_0_0_40 (.A1(n_0_0_83), .A2(n_0_0_82), .ZN(n_0_0_22));
   NOR2_X1 i_0_0_41 (.A1(n_0_0_45), .A2(n_0_0_77), .ZN(n_0_0_20));
   OR2_X1 i_0_0_42 (.A1(n_0_0_77), .A2(n_0_0_76), .ZN(n_0_0_18));
   NAND2_X1 i_0_0_43 (.A1(n_0_0_47), .A2(n_0_0_73), .ZN(n_0_0_16));
   AND2_X1 i_0_0_44 (.A1(n_0_0_73), .A2(n_0_0_72), .ZN(n_0_0_15));
   NOR2_X1 i_0_0_45 (.A1(n_0_0_49), .A2(n_0_0_66), .ZN(n_0_0_13));
   OR2_X1 i_0_0_46 (.A1(n_0_0_66), .A2(n_0_0_65), .ZN(n_0_0_11));
   NAND2_X1 i_0_0_47 (.A1(n_0_0_52), .A2(n_0_0_57), .ZN(n_0_0_9));
   AND2_X1 i_0_0_48 (.A1(n_0_0_57), .A2(n_0_0_56), .ZN(n_0_0_3));
   NAND2_X1 i_0_0_49 (.A1(n_0_0_1), .A2(n_0_0_136), .ZN(negative));
   OAI21_X1 i_0_0_50 (.A(n_0_0_134), .B1(n_0_0_21), .B2(n_0_0_130), .ZN(n_0_0_1));
   INV_X1 i_0_0_51 (.A(n_0_0_2), .ZN(overflow_flag));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_10), .A2(n_0_0_6), .ZN(n_0_0_2));
   NAND3_X1 i_0_0_53 (.A1(n_0_0_19), .A2(n_0_0_134), .A3(n_0_0_129), .ZN(n_0_0_6));
   INV_X1 i_0_0_54 (.A(n_0_0_8), .ZN(carry));
   NAND2_X1 i_0_0_55 (.A1(n_0_0_10), .A2(n_0_0_134), .ZN(n_0_0_8));
   OAI21_X1 i_0_0_56 (.A(n_0_0_136), .B1(n_0_0_21), .B2(n_0_0_130), .ZN(n_0_0_10));
   NAND2_X1 i_0_0_36 (.A1(n_0_0_12), .A2(n_0_0_17), .ZN(result[15]));
   OAI21_X1 i_0_0_37 (.A(n_0_0_14), .B1(n_0_0_21), .B2(n_0_0_130), .ZN(n_0_0_12));
   INV_X1 i_0_0_38 (.A(n_0_0_133), .ZN(n_0_0_14));
   NAND3_X1 i_0_0_39 (.A1(n_0_0_19), .A2(n_0_0_133), .A3(n_0_0_129), .ZN(
      n_0_0_17));
   INV_X1 i_0_0_57 (.A(n_0_0_21), .ZN(n_0_0_19));
   AOI21_X1 i_0_0_58 (.A(n_0_0_127), .B1(n_0_0_24), .B2(n_0_0_124), .ZN(n_0_0_21));
   OAI21_X1 i_0_0_59 (.A(n_0_0_123), .B1(n_0_0_26), .B2(n_0_0_117), .ZN(n_0_0_24));
   AOI21_X1 i_0_0_60 (.A(n_0_0_116), .B1(n_0_0_28), .B2(n_0_0_113), .ZN(n_0_0_26));
   OAI21_X1 i_0_0_61 (.A(n_0_0_112), .B1(n_0_0_31), .B2(n_0_0_107), .ZN(n_0_0_28));
   AOI21_X1 i_0_0_62 (.A(n_0_0_106), .B1(n_0_0_33), .B2(n_0_0_103), .ZN(n_0_0_31));
   OAI21_X1 i_0_0_63 (.A(n_0_0_102), .B1(n_0_0_35), .B2(n_0_0_97), .ZN(n_0_0_33));
   AOI21_X1 i_0_0_64 (.A(n_0_0_96), .B1(n_0_0_38), .B2(n_0_0_93), .ZN(n_0_0_35));
   OAI21_X1 i_0_0_65 (.A(n_0_0_92), .B1(n_0_0_40), .B2(n_0_0_87), .ZN(n_0_0_38));
   AOI21_X1 i_0_0_66 (.A(n_0_0_86), .B1(n_0_0_42), .B2(n_0_0_83), .ZN(n_0_0_40));
   OAI21_X1 i_0_0_67 (.A(n_0_0_82), .B1(n_0_0_45), .B2(n_0_0_77), .ZN(n_0_0_42));
   AOI21_X1 i_0_0_68 (.A(n_0_0_76), .B1(n_0_0_47), .B2(n_0_0_73), .ZN(n_0_0_45));
   OAI21_X1 i_0_0_69 (.A(n_0_0_72), .B1(n_0_0_49), .B2(n_0_0_66), .ZN(n_0_0_47));
   AOI21_X1 i_0_0_70 (.A(n_0_0_65), .B1(n_0_0_52), .B2(n_0_0_57), .ZN(n_0_0_49));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_56), .A2(n_0_0_7), .ZN(n_0_0_52));
   INV_X1 i_0_0_72 (.A(n_0_0_53), .ZN(n_0_0_7));
   NAND2_X1 i_0_0_73 (.A1(n_0_0_5), .A2(n_0_0_55), .ZN(n_0_0_53));
   NAND2_X1 i_0_0_74 (.A1(B[0]), .A2(A[0]), .ZN(n_0_0_55));
   NAND2_X1 i_0_0_75 (.A1(n_0_0_4), .A2(is_subtract), .ZN(n_0_0_5));
   INV_X1 i_0_0_76 (.A(B[0]), .ZN(n_0_0_4));
   NAND3_X1 i_0_0_77 (.A1(n_0_0_62), .A2(A[1]), .A3(n_0_0_59), .ZN(n_0_0_56));
   NAND2_X1 i_0_0_78 (.A1(n_0_0_58), .A2(n_0_0_64), .ZN(n_0_0_57));
   NAND2_X1 i_0_0_79 (.A1(n_0_0_62), .A2(n_0_0_59), .ZN(n_0_0_58));
   NAND2_X1 i_0_0_80 (.A1(B[1]), .A2(is_subtract), .ZN(n_0_0_59));
   NAND2_X1 i_0_0_81 (.A1(n_0_0_63), .A2(n_0_0_121), .ZN(n_0_0_62));
   INV_X1 i_0_0_82 (.A(B[1]), .ZN(n_0_0_63));
   INV_X1 i_0_0_83 (.A(A[1]), .ZN(n_0_0_64));
   AOI21_X1 i_0_0_84 (.A(n_0_0_71), .B1(n_0_0_70), .B2(n_0_0_68), .ZN(n_0_0_65));
   INV_X1 i_0_0_85 (.A(n_0_0_67), .ZN(n_0_0_66));
   NAND3_X1 i_0_0_86 (.A1(n_0_0_70), .A2(n_0_0_68), .A3(n_0_0_71), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_87 (.A1(n_0_0_69), .A2(is_subtract), .ZN(n_0_0_68));
   INV_X1 i_0_0_88 (.A(B[2]), .ZN(n_0_0_69));
   NAND2_X1 i_0_0_89 (.A1(n_0_0_121), .A2(B[2]), .ZN(n_0_0_70));
   INV_X1 i_0_0_90 (.A(A[2]), .ZN(n_0_0_71));
   NAND2_X1 i_0_0_91 (.A1(n_0_0_74), .A2(A[3]), .ZN(n_0_0_72));
   OR2_X1 i_0_0_92 (.A1(n_0_0_74), .A2(A[3]), .ZN(n_0_0_73));
   INV_X1 i_0_0_93 (.A(n_0_0_75), .ZN(n_0_0_74));
   XNOR2_X1 i_0_0_94 (.A(B[3]), .B(is_subtract), .ZN(n_0_0_75));
   NOR2_X1 i_0_0_95 (.A1(n_0_0_79), .A2(n_0_0_81), .ZN(n_0_0_76));
   INV_X1 i_0_0_96 (.A(n_0_0_78), .ZN(n_0_0_77));
   NAND2_X1 i_0_0_97 (.A1(n_0_0_79), .A2(n_0_0_81), .ZN(n_0_0_78));
   INV_X1 i_0_0_98 (.A(n_0_0_80), .ZN(n_0_0_79));
   XNOR2_X1 i_0_0_99 (.A(n_0_0_121), .B(B[4]), .ZN(n_0_0_80));
   INV_X1 i_0_0_100 (.A(A[4]), .ZN(n_0_0_81));
   NAND2_X1 i_0_0_101 (.A1(n_0_0_84), .A2(A[5]), .ZN(n_0_0_82));
   OR2_X1 i_0_0_102 (.A1(n_0_0_84), .A2(A[5]), .ZN(n_0_0_83));
   INV_X1 i_0_0_103 (.A(n_0_0_85), .ZN(n_0_0_84));
   XNOR2_X1 i_0_0_104 (.A(B[5]), .B(is_subtract), .ZN(n_0_0_85));
   NOR2_X1 i_0_0_105 (.A1(n_0_0_89), .A2(n_0_0_91), .ZN(n_0_0_86));
   INV_X1 i_0_0_106 (.A(n_0_0_88), .ZN(n_0_0_87));
   NAND2_X1 i_0_0_107 (.A1(n_0_0_89), .A2(n_0_0_91), .ZN(n_0_0_88));
   INV_X1 i_0_0_108 (.A(n_0_0_90), .ZN(n_0_0_89));
   XNOR2_X1 i_0_0_109 (.A(n_0_0_121), .B(B[6]), .ZN(n_0_0_90));
   INV_X1 i_0_0_110 (.A(A[6]), .ZN(n_0_0_91));
   NAND2_X1 i_0_0_111 (.A1(n_0_0_94), .A2(A[7]), .ZN(n_0_0_92));
   OR2_X1 i_0_0_112 (.A1(n_0_0_94), .A2(A[7]), .ZN(n_0_0_93));
   INV_X1 i_0_0_113 (.A(n_0_0_95), .ZN(n_0_0_94));
   XNOR2_X1 i_0_0_114 (.A(B[7]), .B(is_subtract), .ZN(n_0_0_95));
   NOR2_X1 i_0_0_115 (.A1(n_0_0_99), .A2(n_0_0_101), .ZN(n_0_0_96));
   INV_X1 i_0_0_116 (.A(n_0_0_98), .ZN(n_0_0_97));
   NAND2_X1 i_0_0_117 (.A1(n_0_0_99), .A2(n_0_0_101), .ZN(n_0_0_98));
   INV_X1 i_0_0_118 (.A(n_0_0_100), .ZN(n_0_0_99));
   XNOR2_X1 i_0_0_119 (.A(n_0_0_121), .B(B[8]), .ZN(n_0_0_100));
   INV_X1 i_0_0_120 (.A(A[8]), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_121 (.A1(n_0_0_104), .A2(A[9]), .ZN(n_0_0_102));
   OR2_X1 i_0_0_122 (.A1(n_0_0_104), .A2(A[9]), .ZN(n_0_0_103));
   INV_X1 i_0_0_123 (.A(n_0_0_105), .ZN(n_0_0_104));
   XNOR2_X1 i_0_0_124 (.A(B[9]), .B(is_subtract), .ZN(n_0_0_105));
   NOR2_X1 i_0_0_125 (.A1(n_0_0_109), .A2(n_0_0_111), .ZN(n_0_0_106));
   INV_X1 i_0_0_126 (.A(n_0_0_108), .ZN(n_0_0_107));
   NAND2_X1 i_0_0_127 (.A1(n_0_0_109), .A2(n_0_0_111), .ZN(n_0_0_108));
   INV_X1 i_0_0_128 (.A(n_0_0_110), .ZN(n_0_0_109));
   XNOR2_X1 i_0_0_129 (.A(n_0_0_121), .B(B[10]), .ZN(n_0_0_110));
   INV_X1 i_0_0_130 (.A(A[10]), .ZN(n_0_0_111));
   NAND2_X1 i_0_0_131 (.A1(n_0_0_114), .A2(A[11]), .ZN(n_0_0_112));
   OR2_X1 i_0_0_132 (.A1(n_0_0_114), .A2(A[11]), .ZN(n_0_0_113));
   INV_X1 i_0_0_133 (.A(n_0_0_115), .ZN(n_0_0_114));
   XNOR2_X1 i_0_0_134 (.A(B[11]), .B(is_subtract), .ZN(n_0_0_115));
   NOR2_X1 i_0_0_135 (.A1(n_0_0_119), .A2(n_0_0_122), .ZN(n_0_0_116));
   INV_X1 i_0_0_136 (.A(n_0_0_118), .ZN(n_0_0_117));
   NAND2_X1 i_0_0_137 (.A1(n_0_0_119), .A2(n_0_0_122), .ZN(n_0_0_118));
   INV_X1 i_0_0_138 (.A(n_0_0_120), .ZN(n_0_0_119));
   XNOR2_X1 i_0_0_139 (.A(n_0_0_121), .B(B[12]), .ZN(n_0_0_120));
   INV_X1 i_0_0_140 (.A(is_subtract), .ZN(n_0_0_121));
   INV_X1 i_0_0_141 (.A(A[12]), .ZN(n_0_0_122));
   NAND2_X1 i_0_0_142 (.A1(n_0_0_125), .A2(A[13]), .ZN(n_0_0_123));
   OR2_X1 i_0_0_143 (.A1(n_0_0_125), .A2(A[13]), .ZN(n_0_0_124));
   INV_X1 i_0_0_144 (.A(n_0_0_126), .ZN(n_0_0_125));
   XNOR2_X1 i_0_0_145 (.A(B[13]), .B(is_subtract), .ZN(n_0_0_126));
   INV_X1 i_0_0_146 (.A(n_0_0_128), .ZN(n_0_0_127));
   NAND2_X1 i_0_0_147 (.A1(n_0_0_131), .A2(A[14]), .ZN(n_0_0_128));
   INV_X1 i_0_0_148 (.A(n_0_0_130), .ZN(n_0_0_129));
   NOR2_X1 i_0_0_149 (.A1(n_0_0_131), .A2(A[14]), .ZN(n_0_0_130));
   INV_X1 i_0_0_150 (.A(n_0_0_132), .ZN(n_0_0_131));
   XNOR2_X1 i_0_0_151 (.A(B[14]), .B(is_subtract), .ZN(n_0_0_132));
   NAND2_X1 i_0_0_152 (.A1(n_0_0_134), .A2(n_0_0_136), .ZN(n_0_0_133));
   INV_X1 i_0_0_153 (.A(n_0_0_135), .ZN(n_0_0_134));
   NOR2_X1 i_0_0_154 (.A1(n_0_0_0), .A2(A[15]), .ZN(n_0_0_135));
   NAND2_X1 i_0_0_155 (.A1(n_0_0_0), .A2(A[15]), .ZN(n_0_0_136));
endmodule
