/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Apr 24 00:11:39 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 757929726 */

module RAM_after(clk, rst, we1, addr1, addr2, data1, data2);
   input clk;
   input rst;
   input we1;
   input [3:0]addr1;
   input [3:0]addr2;
   inout [31:0]data1;
   output [31:0]data2;

   wire n_32_0;
   wire [31:0]\MEM[15] ;
   wire n_32_1;
   wire [31:0]\MEM[14] ;
   wire n_32_2;
   wire [31:0]\MEM[13] ;
   wire n_32_3;
   wire [31:0]\MEM[12] ;
   wire n_32_4;
   wire [31:0]\MEM[11] ;
   wire n_32_5;
   wire [31:0]\MEM[10] ;
   wire n_32_6;
   wire [31:0]\MEM[9] ;
   wire n_32_7;
   wire [31:0]\MEM[8] ;
   wire n_32_8;
   wire [31:0]\MEM[7] ;
   wire n_32_9;
   wire [31:0]\MEM[6] ;
   wire n_32_10;
   wire [31:0]\MEM[5] ;
   wire n_32_11;
   wire [31:0]\MEM[4] ;
   wire n_32_12;
   wire [31:0]\MEM[3] ;
   wire n_32_13;
   wire [31:0]\MEM[2] ;
   wire n_32_14;
   wire [31:0]\MEM[1] ;
   wire n_32_15;
   wire [31:0]\MEM[0] ;
   wire n_32_0_0;
   wire n_32_0_1;
   wire n_32_0_2;
   wire n_32_0_3;
   wire n_32_0_4;
   wire n_32_0_5;
   wire n_32_0_6;
   wire n_32_0_7;
   wire n_32_0_8;
   wire n_32_0_9;
   wire n_32_0_10;
   wire n_32_0_11;
   wire n_32_0_12;
   wire n_32_0_13;
   wire n_32_0_14;
   wire n_32_0_15;
   wire n_32_0_16;
   wire n_32_0_17;
   wire n_32_0_18;
   wire n_32_0_19;
   wire n_32_0_20;
   wire n_32_0_21;
   wire n_32_0_22;
   wire n_32_0_23;
   wire n_32_0_24;
   wire n_32_0_25;
   wire n_32_0_26;
   wire n_32_0_27;
   wire n_32_0_28;
   wire n_32_0_29;
   wire n_32_0_30;
   wire n_32_0_31;
   wire n_32_0_32;
   wire n_32_0_33;
   wire n_32_0_34;
   wire [31:0]MEM;
   wire n_32_0_35;
   wire n_32_0_36;
   wire n_32_16;
   wire n_32_0_37;
   wire n_32_0_38;
   wire n_32_0_39;
   wire n_32_0_40;
   wire n_32_0_41;
   wire n_32_0_42;
   wire n_32_0_43;
   wire n_32_0_44;
   wire n_32_0_45;
   wire n_32_0_46;
   wire n_32_17;
   wire n_32_0_47;
   wire n_32_0_48;
   wire n_32_0_49;
   wire n_32_0_50;
   wire n_32_0_51;
   wire n_32_0_52;
   wire n_32_0_53;
   wire n_32_0_54;
   wire n_32_0_55;
   wire n_32_0_56;
   wire n_32_18;
   wire n_32_0_57;
   wire n_32_0_58;
   wire n_32_0_59;
   wire n_32_0_60;
   wire n_32_0_61;
   wire n_32_0_62;
   wire n_32_0_63;
   wire n_32_0_64;
   wire n_32_0_65;
   wire n_32_0_66;
   wire n_32_19;
   wire n_32_0_67;
   wire n_32_0_68;
   wire n_32_0_69;
   wire n_32_0_70;
   wire n_32_0_71;
   wire n_32_0_72;
   wire n_32_0_73;
   wire n_32_0_74;
   wire n_32_0_75;
   wire n_32_0_76;
   wire n_32_20;
   wire n_32_0_77;
   wire n_32_0_78;
   wire n_32_0_79;
   wire n_32_0_80;
   wire n_32_0_81;
   wire n_32_0_82;
   wire n_32_0_83;
   wire n_32_0_84;
   wire n_32_0_85;
   wire n_32_0_86;
   wire n_32_21;
   wire n_32_0_87;
   wire n_32_0_88;
   wire n_32_0_89;
   wire n_32_0_90;
   wire n_32_0_91;
   wire n_32_0_92;
   wire n_32_0_93;
   wire n_32_0_94;
   wire n_32_0_95;
   wire n_32_0_96;
   wire n_32_22;
   wire n_32_0_97;
   wire n_32_0_98;
   wire n_32_0_99;
   wire n_32_0_100;
   wire n_32_0_101;
   wire n_32_0_102;
   wire n_32_0_103;
   wire n_32_0_104;
   wire n_32_0_105;
   wire n_32_0_106;
   wire n_32_23;
   wire n_32_0_107;
   wire n_32_0_108;
   wire n_32_0_109;
   wire n_32_0_110;
   wire n_32_0_111;
   wire n_32_0_112;
   wire n_32_0_113;
   wire n_32_0_114;
   wire n_32_0_115;
   wire n_32_0_116;
   wire n_32_24;
   wire n_32_0_117;
   wire n_32_0_118;
   wire n_32_0_119;
   wire n_32_0_120;
   wire n_32_0_121;
   wire n_32_0_122;
   wire n_32_0_123;
   wire n_32_0_124;
   wire n_32_0_125;
   wire n_32_0_126;
   wire n_32_25;
   wire n_32_0_127;
   wire n_32_0_128;
   wire n_32_0_129;
   wire n_32_0_130;
   wire n_32_0_131;
   wire n_32_0_132;
   wire n_32_0_133;
   wire n_32_0_134;
   wire n_32_0_135;
   wire n_32_0_136;
   wire n_32_26;
   wire n_32_0_137;
   wire n_32_0_138;
   wire n_32_0_139;
   wire n_32_0_140;
   wire n_32_0_141;
   wire n_32_0_142;
   wire n_32_0_143;
   wire n_32_0_144;
   wire n_32_0_145;
   wire n_32_0_146;
   wire n_32_27;
   wire n_32_0_147;
   wire n_32_0_148;
   wire n_32_0_149;
   wire n_32_0_150;
   wire n_32_0_151;
   wire n_32_0_152;
   wire n_32_0_153;
   wire n_32_0_154;
   wire n_32_0_155;
   wire n_32_0_156;
   wire n_32_28;
   wire n_32_0_157;
   wire n_32_0_158;
   wire n_32_0_159;
   wire n_32_0_160;
   wire n_32_0_161;
   wire n_32_0_162;
   wire n_32_0_163;
   wire n_32_0_164;
   wire n_32_0_165;
   wire n_32_0_166;
   wire n_32_29;
   wire n_32_0_167;
   wire n_32_0_168;
   wire n_32_0_169;
   wire n_32_0_170;
   wire n_32_0_171;
   wire n_32_0_172;
   wire n_32_0_173;
   wire n_32_0_174;
   wire n_32_0_175;
   wire n_32_0_176;
   wire n_32_30;
   wire n_32_0_177;
   wire n_32_0_178;
   wire n_32_0_179;
   wire n_32_0_180;
   wire n_32_0_181;
   wire n_32_0_182;
   wire n_32_0_183;
   wire n_32_0_184;
   wire n_32_0_185;
   wire n_32_0_186;
   wire n_32_31;
   wire n_32_0_187;
   wire n_32_0_188;
   wire n_32_0_189;
   wire n_32_0_190;
   wire n_32_0_191;
   wire n_32_0_192;
   wire n_32_0_193;
   wire n_32_0_194;
   wire n_32_0_195;
   wire n_32_0_196;
   wire n_32_32;
   wire n_32_0_197;
   wire n_32_0_198;
   wire n_32_0_199;
   wire n_32_0_200;
   wire n_32_0_201;
   wire n_32_0_202;
   wire n_32_0_203;
   wire n_32_0_204;
   wire n_32_0_205;
   wire n_32_0_206;
   wire n_32_33;
   wire n_32_0_207;
   wire n_32_0_208;
   wire n_32_0_209;
   wire n_32_0_210;
   wire n_32_0_211;
   wire n_32_0_212;
   wire n_32_0_213;
   wire n_32_0_214;
   wire n_32_0_215;
   wire n_32_0_216;
   wire n_32_34;
   wire n_32_0_217;
   wire n_32_0_218;
   wire n_32_0_219;
   wire n_32_0_220;
   wire n_32_0_221;
   wire n_32_0_222;
   wire n_32_0_223;
   wire n_32_0_224;
   wire n_32_0_225;
   wire n_32_0_226;
   wire n_32_35;
   wire n_32_0_227;
   wire n_32_0_228;
   wire n_32_0_229;
   wire n_32_0_230;
   wire n_32_0_231;
   wire n_32_0_232;
   wire n_32_0_233;
   wire n_32_0_234;
   wire n_32_0_235;
   wire n_32_0_236;
   wire n_32_36;
   wire n_32_0_237;
   wire n_32_0_238;
   wire n_32_0_239;
   wire n_32_0_240;
   wire n_32_0_241;
   wire n_32_0_242;
   wire n_32_0_243;
   wire n_32_0_244;
   wire n_32_0_245;
   wire n_32_0_246;
   wire n_32_37;
   wire n_32_0_247;
   wire n_32_0_248;
   wire n_32_0_249;
   wire n_32_0_250;
   wire n_32_0_251;
   wire n_32_0_252;
   wire n_32_0_253;
   wire n_32_0_254;
   wire n_32_0_255;
   wire n_32_0_256;
   wire n_32_38;
   wire n_32_0_257;
   wire n_32_0_258;
   wire n_32_0_259;
   wire n_32_0_260;
   wire n_32_0_261;
   wire n_32_0_262;
   wire n_32_0_263;
   wire n_32_0_264;
   wire n_32_0_265;
   wire n_32_0_266;
   wire n_32_39;
   wire n_32_0_267;
   wire n_32_0_268;
   wire n_32_0_269;
   wire n_32_0_270;
   wire n_32_0_271;
   wire n_32_0_272;
   wire n_32_0_273;
   wire n_32_0_274;
   wire n_32_0_275;
   wire n_32_0_276;
   wire n_32_40;
   wire n_32_0_277;
   wire n_32_0_278;
   wire n_32_0_279;
   wire n_32_0_280;
   wire n_32_0_281;
   wire n_32_0_282;
   wire n_32_0_283;
   wire n_32_0_284;
   wire n_32_0_285;
   wire n_32_0_286;
   wire n_32_41;
   wire n_32_0_287;
   wire n_32_0_288;
   wire n_32_0_289;
   wire n_32_0_290;
   wire n_32_0_291;
   wire n_32_0_292;
   wire n_32_0_293;
   wire n_32_0_294;
   wire n_32_0_295;
   wire n_32_0_296;
   wire n_32_42;
   wire n_32_0_297;
   wire n_32_0_298;
   wire n_32_0_299;
   wire n_32_0_300;
   wire n_32_0_301;
   wire n_32_0_302;
   wire n_32_0_303;
   wire n_32_0_304;
   wire n_32_0_305;
   wire n_32_0_306;
   wire n_32_43;
   wire n_32_0_307;
   wire n_32_0_308;
   wire n_32_0_309;
   wire n_32_0_310;
   wire n_32_0_311;
   wire n_32_0_312;
   wire n_32_0_313;
   wire n_32_0_314;
   wire n_32_0_315;
   wire n_32_0_316;
   wire n_32_44;
   wire n_32_0_317;
   wire n_32_0_318;
   wire n_32_0_319;
   wire n_32_0_320;
   wire n_32_0_321;
   wire n_32_0_322;
   wire n_32_0_323;
   wire n_32_0_324;
   wire n_32_0_325;
   wire n_32_0_326;
   wire n_32_45;
   wire n_32_0_327;
   wire n_32_0_328;
   wire n_32_0_329;
   wire n_32_0_330;
   wire n_32_0_331;
   wire n_32_0_332;
   wire n_32_0_333;
   wire n_32_0_334;
   wire n_32_0_335;
   wire n_32_0_336;
   wire n_32_46;
   wire n_32_0_337;
   wire n_32_0_338;
   wire n_32_0_339;
   wire n_32_0_340;
   wire n_32_0_341;
   wire n_32_0_342;
   wire n_32_0_343;
   wire n_32_0_344;
   wire n_32_0_345;
   wire n_32_0_346;
   wire n_32_0_347;
   wire n_32_0_348;
   wire n_32_47;
   wire n_32_48;
   wire n_32_49;
   wire n_32_50;
   wire n_32_51;
   wire n_32_52;
   wire n_32_53;
   wire n_32_54;
   wire n_32_55;
   wire n_32_56;
   wire n_32_57;
   wire n_32_58;
   wire n_32_59;
   wire n_32_60;
   wire n_32_61;
   wire n_32_62;
   wire n_32_63;
   wire n_32_0_349;
   wire n_32_0_350;
   wire n_32_0_351;
   wire n_32_0_352;
   wire n_32_0_353;
   wire n_32_0_354;
   wire n_32_0_355;
   wire n_32_0_356;
   wire n_32_0_357;
   wire n_32_0_358;
   wire n_32_0_359;
   wire n_32_0_360;
   wire n_32_0_361;
   wire n_32_0_362;
   wire n_32_0_363;
   wire n_32_0_364;
   wire n_32_0_365;
   wire n_32_0_366;
   wire n_32_0_367;
   wire n_32_0_368;
   wire n_32_0_369;
   wire n_32_0_370;
   wire n_32_0_371;
   wire n_32_0_372;
   wire n_32_0_373;
   wire n_32_0_374;
   wire n_32_0_375;
   wire n_32_0_376;
   wire n_32_0_377;
   wire n_32_0_378;
   wire n_32_0_379;
   wire n_32_0_380;
   wire n_32_0_381;
   wire n_32_0_382;
   wire n_32_0_383;
   wire n_32_0_384;
   wire n_32_0_385;
   wire n_32_0_386;
   wire n_32_0_387;
   wire n_32_0_388;
   wire n_32_0_389;
   wire n_32_0_390;
   wire n_32_0_391;
   wire n_32_0_392;
   wire n_32_0_393;
   wire n_32_0_394;
   wire n_32_0_395;
   wire n_32_0_396;
   wire n_32_0_397;
   wire n_32_0_398;
   wire n_32_0_399;
   wire n_32_0_400;
   wire n_32_0_401;
   wire n_32_0_402;
   wire n_32_0_403;
   wire n_32_0_404;
   wire n_32_0_405;
   wire n_32_0_406;
   wire n_32_0_407;
   wire n_32_0_408;
   wire n_32_0_409;
   wire n_32_0_410;
   wire n_32_0_411;
   wire n_32_0_412;
   wire n_32_0_413;
   wire n_32_0_414;
   wire n_32_0_415;
   wire n_32_0_416;
   wire n_32_0_417;
   wire n_32_0_418;
   wire n_32_0_419;
   wire n_32_0_420;
   wire n_32_0_421;
   wire n_32_0_422;
   wire n_32_0_423;
   wire n_32_0_424;
   wire n_32_0_425;
   wire n_32_0_426;
   wire n_32_0_427;
   wire n_32_0_428;
   wire n_32_0_429;
   wire n_32_0_430;
   wire n_32_0_431;
   wire n_32_0_432;
   wire n_32_0_433;
   wire n_32_0_434;
   wire n_32_0_435;
   wire n_32_0_436;
   wire n_32_0_437;
   wire n_32_0_438;
   wire n_32_0_439;
   wire n_32_0_440;
   wire n_32_0_441;
   wire n_32_0_442;
   wire n_32_0_443;
   wire n_32_0_444;
   wire n_32_0_445;
   wire n_32_0_446;
   wire n_32_0_447;
   wire n_32_0_448;
   wire n_32_0_449;
   wire n_32_0_450;
   wire n_32_0_451;
   wire n_32_0_452;
   wire n_32_0_453;
   wire n_32_0_454;
   wire n_32_0_455;
   wire n_32_0_456;
   wire n_32_0_457;
   wire n_32_0_458;
   wire n_32_0_459;
   wire n_32_0_460;
   wire n_32_0_461;
   wire n_32_0_462;
   wire n_32_0_463;
   wire n_32_0_464;
   wire n_32_0_465;
   wire n_32_0_466;
   wire n_32_0_467;
   wire n_32_0_468;
   wire n_32_0_469;
   wire n_32_0_470;
   wire n_32_0_471;
   wire n_32_0_472;
   wire n_32_0_473;
   wire n_32_0_474;
   wire n_32_0_475;
   wire n_32_0_476;
   wire n_32_0_477;
   wire n_32_0_478;
   wire n_32_0_479;
   wire n_32_0_480;
   wire n_32_0_481;
   wire n_32_0_482;
   wire n_32_0_483;
   wire n_32_0_484;
   wire n_32_0_485;
   wire n_32_0_486;
   wire n_32_0_487;
   wire n_32_0_488;
   wire n_32_0_489;
   wire n_32_0_490;
   wire n_32_0_491;
   wire n_32_0_492;
   wire n_32_0_493;
   wire n_32_0_494;
   wire n_32_0_495;
   wire n_32_0_496;
   wire n_32_0_497;
   wire n_32_0_498;
   wire n_32_0_499;
   wire n_32_0_500;
   wire n_32_0_501;
   wire n_32_0_502;
   wire n_32_0_503;
   wire n_32_0_504;
   wire n_32_0_505;
   wire n_32_0_506;
   wire n_32_0_507;
   wire n_32_0_508;
   wire n_32_0_509;
   wire n_32_0_510;
   wire n_32_0_511;
   wire n_32_0_512;
   wire n_32_0_513;
   wire n_32_0_514;
   wire n_32_0_515;
   wire n_32_0_516;
   wire n_32_0_517;
   wire n_32_0_518;
   wire n_32_0_519;
   wire n_32_0_520;
   wire n_32_0_521;
   wire n_32_0_522;
   wire n_32_0_523;
   wire n_32_0_524;
   wire n_32_0_525;
   wire n_32_0_526;
   wire n_32_0_527;
   wire n_32_0_528;
   wire n_32_0_529;
   wire n_32_0_530;
   wire n_32_0_531;
   wire n_32_0_532;
   wire n_32_0_533;
   wire n_32_0_534;
   wire n_32_0_535;
   wire n_32_0_536;
   wire n_32_0_537;
   wire n_32_0_538;
   wire n_32_0_539;
   wire n_32_0_540;
   wire n_32_0_541;
   wire n_32_0_542;
   wire n_32_0_543;
   wire n_32_0_544;
   wire n_32_0_545;
   wire n_32_0_546;
   wire n_32_0_547;
   wire n_32_0_548;
   wire n_32_0_549;
   wire n_32_0_550;
   wire n_32_0_551;
   wire n_32_0_552;
   wire n_32_0_553;
   wire n_32_0_554;
   wire n_32_0_555;
   wire n_32_0_556;
   wire n_32_0_557;
   wire n_32_0_558;
   wire n_32_0_559;
   wire n_32_0_560;
   wire n_32_0_561;
   wire n_32_0_562;
   wire n_32_0_563;
   wire n_32_0_564;
   wire n_32_0_565;
   wire n_32_0_566;
   wire n_32_0_567;
   wire n_32_0_568;
   wire n_32_0_569;
   wire n_32_0_570;
   wire n_32_0_571;
   wire n_32_0_572;
   wire n_32_0_573;
   wire n_32_0_574;
   wire n_32_0_575;
   wire n_32_0_576;
   wire n_32_0_577;
   wire n_32_0_578;
   wire n_32_0_579;
   wire n_32_0_580;
   wire n_32_0_581;
   wire n_32_0_582;
   wire n_32_0_583;
   wire n_32_0_584;
   wire n_32_0_585;
   wire n_32_0_586;
   wire n_32_0_587;
   wire n_32_0_588;
   wire n_32_0_589;
   wire n_32_0_590;
   wire n_32_0_591;
   wire n_32_0_592;
   wire n_32_0_593;
   wire n_32_0_594;
   wire n_32_0_595;
   wire n_32_0_596;
   wire n_32_0_597;
   wire n_32_0_598;
   wire n_32_0_599;
   wire n_32_0_600;
   wire n_32_0_601;
   wire n_32_0_602;
   wire n_32_0_603;
   wire n_32_0_604;
   wire n_32_0_605;
   wire n_32_0_606;
   wire n_32_0_607;
   wire n_32_0_608;
   wire n_32_0_609;
   wire n_32_0_610;
   wire n_32_0_611;
   wire n_32_0_612;
   wire n_32_0_613;
   wire n_32_0_614;
   wire n_32_0_615;
   wire n_32_0_616;
   wire n_32_0_617;
   wire n_32_0_618;
   wire n_32_0_619;
   wire n_32_0_620;
   wire n_32_0_621;
   wire n_32_0_622;
   wire n_32_0_623;
   wire n_32_0_624;
   wire n_32_0_625;
   wire n_32_0_626;
   wire n_32_0_627;
   wire n_32_0_628;
   wire n_32_0_629;
   wire n_32_0_630;
   wire n_32_0_631;
   wire n_32_0_632;
   wire n_32_0_633;
   wire n_32_0_634;
   wire n_32_0_635;
   wire n_32_0_636;
   wire n_32_0_637;
   wire n_32_0_638;
   wire n_32_0_639;
   wire n_32_0_640;
   wire n_32_0_641;
   wire n_32_0_642;
   wire n_32_0_643;
   wire n_32_0_644;
   wire n_32_0_645;
   wire n_32_0_646;
   wire n_32_0_647;
   wire n_32_0_648;
   wire n_32_0_649;
   wire n_32_0_650;
   wire n_32_0_651;
   wire n_32_0_652;
   wire n_32_0_653;
   wire n_32_0_654;
   wire n_32_0_655;
   wire n_32_0_656;
   wire n_32_0_657;
   wire n_32_0_658;
   wire n_32_0_659;
   wire n_32_0_660;
   wire n_32_0_661;
   wire n_32_0_662;
   wire n_32_0_663;
   wire n_32_0_664;
   wire n_32_0_665;
   wire n_32_0_666;
   wire n_32_0_667;

   TBUF_X1 i_0 (.A(MEM[0]), .EN(we1), .Z(data1[0]));
   TBUF_X1 i_1 (.A(MEM[1]), .EN(we1), .Z(data1[1]));
   TBUF_X1 i_2 (.A(MEM[2]), .EN(we1), .Z(data1[2]));
   TBUF_X1 i_3 (.A(MEM[3]), .EN(we1), .Z(data1[3]));
   TBUF_X1 i_4 (.A(MEM[4]), .EN(we1), .Z(data1[4]));
   TBUF_X1 i_5 (.A(MEM[5]), .EN(we1), .Z(data1[5]));
   TBUF_X1 i_6 (.A(MEM[6]), .EN(we1), .Z(data1[6]));
   TBUF_X1 i_7 (.A(MEM[7]), .EN(we1), .Z(data1[7]));
   TBUF_X1 i_8 (.A(MEM[8]), .EN(we1), .Z(data1[8]));
   TBUF_X1 i_9 (.A(MEM[9]), .EN(we1), .Z(data1[9]));
   TBUF_X1 i_10 (.A(MEM[10]), .EN(we1), .Z(data1[10]));
   TBUF_X1 i_11 (.A(MEM[11]), .EN(we1), .Z(data1[11]));
   TBUF_X1 i_12 (.A(MEM[12]), .EN(we1), .Z(data1[12]));
   TBUF_X1 i_13 (.A(MEM[13]), .EN(we1), .Z(data1[13]));
   TBUF_X1 i_14 (.A(MEM[14]), .EN(we1), .Z(data1[14]));
   TBUF_X1 i_15 (.A(MEM[15]), .EN(we1), .Z(data1[15]));
   TBUF_X1 i_16 (.A(MEM[16]), .EN(we1), .Z(data1[16]));
   TBUF_X1 i_17 (.A(MEM[17]), .EN(we1), .Z(data1[17]));
   TBUF_X1 i_18 (.A(MEM[18]), .EN(we1), .Z(data1[18]));
   TBUF_X1 i_19 (.A(MEM[19]), .EN(we1), .Z(data1[19]));
   TBUF_X1 i_20 (.A(MEM[20]), .EN(we1), .Z(data1[20]));
   TBUF_X1 i_21 (.A(MEM[21]), .EN(we1), .Z(data1[21]));
   TBUF_X1 i_22 (.A(MEM[22]), .EN(we1), .Z(data1[22]));
   TBUF_X1 i_23 (.A(MEM[23]), .EN(we1), .Z(data1[23]));
   TBUF_X1 i_24 (.A(MEM[24]), .EN(we1), .Z(data1[24]));
   TBUF_X1 i_25 (.A(MEM[25]), .EN(we1), .Z(data1[25]));
   TBUF_X1 i_26 (.A(MEM[26]), .EN(we1), .Z(data1[26]));
   TBUF_X1 i_27 (.A(MEM[27]), .EN(we1), .Z(data1[27]));
   TBUF_X1 i_28 (.A(MEM[28]), .EN(we1), .Z(data1[28]));
   TBUF_X1 i_29 (.A(MEM[29]), .EN(we1), .Z(data1[29]));
   TBUF_X1 i_30 (.A(MEM[30]), .EN(we1), .Z(data1[30]));
   TBUF_X1 i_31 (.A(MEM[31]), .EN(we1), .Z(data1[31]));
   CLKGATETST_X1 \clk_gate_MEM_reg[15]_reg  (.CK(clk), .E(n_32_63), .SE(1'b0), 
      .GCK(n_32_0));
   DFF_X1 \MEM_reg[15][31]  (.D(n_32_47), .CK(n_32_0), .Q(\MEM[15] [31]), .QN());
   DFF_X1 \MEM_reg[15][30]  (.D(n_32_46), .CK(n_32_0), .Q(\MEM[15] [30]), .QN());
   DFF_X1 \MEM_reg[15][29]  (.D(n_32_45), .CK(n_32_0), .Q(\MEM[15] [29]), .QN());
   DFF_X1 \MEM_reg[15][28]  (.D(n_32_44), .CK(n_32_0), .Q(\MEM[15] [28]), .QN());
   DFF_X1 \MEM_reg[15][27]  (.D(n_32_43), .CK(n_32_0), .Q(\MEM[15] [27]), .QN());
   DFF_X1 \MEM_reg[15][26]  (.D(n_32_42), .CK(n_32_0), .Q(\MEM[15] [26]), .QN());
   DFF_X1 \MEM_reg[15][25]  (.D(n_32_41), .CK(n_32_0), .Q(\MEM[15] [25]), .QN());
   DFF_X1 \MEM_reg[15][24]  (.D(n_32_40), .CK(n_32_0), .Q(\MEM[15] [24]), .QN());
   DFF_X1 \MEM_reg[15][23]  (.D(n_32_39), .CK(n_32_0), .Q(\MEM[15] [23]), .QN());
   DFF_X1 \MEM_reg[15][22]  (.D(n_32_38), .CK(n_32_0), .Q(\MEM[15] [22]), .QN());
   DFF_X1 \MEM_reg[15][21]  (.D(n_32_37), .CK(n_32_0), .Q(\MEM[15] [21]), .QN());
   DFF_X1 \MEM_reg[15][20]  (.D(n_32_36), .CK(n_32_0), .Q(\MEM[15] [20]), .QN());
   DFF_X1 \MEM_reg[15][19]  (.D(n_32_35), .CK(n_32_0), .Q(\MEM[15] [19]), .QN());
   DFF_X1 \MEM_reg[15][18]  (.D(n_32_34), .CK(n_32_0), .Q(\MEM[15] [18]), .QN());
   DFF_X1 \MEM_reg[15][17]  (.D(n_32_33), .CK(n_32_0), .Q(\MEM[15] [17]), .QN());
   DFF_X1 \MEM_reg[15][16]  (.D(n_32_32), .CK(n_32_0), .Q(\MEM[15] [16]), .QN());
   DFF_X1 \MEM_reg[15][15]  (.D(n_32_31), .CK(n_32_0), .Q(\MEM[15] [15]), .QN());
   DFF_X1 \MEM_reg[15][14]  (.D(n_32_30), .CK(n_32_0), .Q(\MEM[15] [14]), .QN());
   DFF_X1 \MEM_reg[15][13]  (.D(n_32_29), .CK(n_32_0), .Q(\MEM[15] [13]), .QN());
   DFF_X1 \MEM_reg[15][12]  (.D(n_32_28), .CK(n_32_0), .Q(\MEM[15] [12]), .QN());
   DFF_X1 \MEM_reg[15][11]  (.D(n_32_27), .CK(n_32_0), .Q(\MEM[15] [11]), .QN());
   DFF_X1 \MEM_reg[15][10]  (.D(n_32_26), .CK(n_32_0), .Q(\MEM[15] [10]), .QN());
   DFF_X1 \MEM_reg[15][9]  (.D(n_32_25), .CK(n_32_0), .Q(\MEM[15] [9]), .QN());
   DFF_X1 \MEM_reg[15][8]  (.D(n_32_24), .CK(n_32_0), .Q(\MEM[15] [8]), .QN());
   DFF_X1 \MEM_reg[15][7]  (.D(n_32_23), .CK(n_32_0), .Q(\MEM[15] [7]), .QN());
   DFF_X1 \MEM_reg[15][6]  (.D(n_32_22), .CK(n_32_0), .Q(\MEM[15] [6]), .QN());
   DFF_X1 \MEM_reg[15][5]  (.D(n_32_21), .CK(n_32_0), .Q(\MEM[15] [5]), .QN());
   DFF_X1 \MEM_reg[15][4]  (.D(n_32_20), .CK(n_32_0), .Q(\MEM[15] [4]), .QN());
   DFF_X1 \MEM_reg[15][3]  (.D(n_32_19), .CK(n_32_0), .Q(\MEM[15] [3]), .QN());
   DFF_X1 \MEM_reg[15][2]  (.D(n_32_18), .CK(n_32_0), .Q(\MEM[15] [2]), .QN());
   DFF_X1 \MEM_reg[15][1]  (.D(n_32_17), .CK(n_32_0), .Q(\MEM[15] [1]), .QN());
   DFF_X1 \MEM_reg[15][0]  (.D(n_32_16), .CK(n_32_0), .Q(\MEM[15] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[14]_reg  (.CK(clk), .E(n_32_62), .SE(1'b0), 
      .GCK(n_32_1));
   DFF_X1 \MEM_reg[14][31]  (.D(n_32_47), .CK(n_32_1), .Q(\MEM[14] [31]), .QN());
   DFF_X1 \MEM_reg[14][30]  (.D(n_32_46), .CK(n_32_1), .Q(\MEM[14] [30]), .QN());
   DFF_X1 \MEM_reg[14][29]  (.D(n_32_45), .CK(n_32_1), .Q(\MEM[14] [29]), .QN());
   DFF_X1 \MEM_reg[14][28]  (.D(n_32_44), .CK(n_32_1), .Q(\MEM[14] [28]), .QN());
   DFF_X1 \MEM_reg[14][27]  (.D(n_32_43), .CK(n_32_1), .Q(\MEM[14] [27]), .QN());
   DFF_X1 \MEM_reg[14][26]  (.D(n_32_42), .CK(n_32_1), .Q(\MEM[14] [26]), .QN());
   DFF_X1 \MEM_reg[14][25]  (.D(n_32_41), .CK(n_32_1), .Q(\MEM[14] [25]), .QN());
   DFF_X1 \MEM_reg[14][24]  (.D(n_32_40), .CK(n_32_1), .Q(\MEM[14] [24]), .QN());
   DFF_X1 \MEM_reg[14][23]  (.D(n_32_39), .CK(n_32_1), .Q(\MEM[14] [23]), .QN());
   DFF_X1 \MEM_reg[14][22]  (.D(n_32_38), .CK(n_32_1), .Q(\MEM[14] [22]), .QN());
   DFF_X1 \MEM_reg[14][21]  (.D(n_32_37), .CK(n_32_1), .Q(\MEM[14] [21]), .QN());
   DFF_X1 \MEM_reg[14][20]  (.D(n_32_36), .CK(n_32_1), .Q(\MEM[14] [20]), .QN());
   DFF_X1 \MEM_reg[14][19]  (.D(n_32_35), .CK(n_32_1), .Q(\MEM[14] [19]), .QN());
   DFF_X1 \MEM_reg[14][18]  (.D(n_32_34), .CK(n_32_1), .Q(\MEM[14] [18]), .QN());
   DFF_X1 \MEM_reg[14][17]  (.D(n_32_33), .CK(n_32_1), .Q(\MEM[14] [17]), .QN());
   DFF_X1 \MEM_reg[14][16]  (.D(n_32_32), .CK(n_32_1), .Q(\MEM[14] [16]), .QN());
   DFF_X1 \MEM_reg[14][15]  (.D(n_32_31), .CK(n_32_1), .Q(\MEM[14] [15]), .QN());
   DFF_X1 \MEM_reg[14][14]  (.D(n_32_30), .CK(n_32_1), .Q(\MEM[14] [14]), .QN());
   DFF_X1 \MEM_reg[14][13]  (.D(n_32_29), .CK(n_32_1), .Q(\MEM[14] [13]), .QN());
   DFF_X1 \MEM_reg[14][12]  (.D(n_32_28), .CK(n_32_1), .Q(\MEM[14] [12]), .QN());
   DFF_X1 \MEM_reg[14][11]  (.D(n_32_27), .CK(n_32_1), .Q(\MEM[14] [11]), .QN());
   DFF_X1 \MEM_reg[14][10]  (.D(n_32_26), .CK(n_32_1), .Q(\MEM[14] [10]), .QN());
   DFF_X1 \MEM_reg[14][9]  (.D(n_32_25), .CK(n_32_1), .Q(\MEM[14] [9]), .QN());
   DFF_X1 \MEM_reg[14][8]  (.D(n_32_24), .CK(n_32_1), .Q(\MEM[14] [8]), .QN());
   DFF_X1 \MEM_reg[14][7]  (.D(n_32_23), .CK(n_32_1), .Q(\MEM[14] [7]), .QN());
   DFF_X1 \MEM_reg[14][6]  (.D(n_32_22), .CK(n_32_1), .Q(\MEM[14] [6]), .QN());
   DFF_X1 \MEM_reg[14][5]  (.D(n_32_21), .CK(n_32_1), .Q(\MEM[14] [5]), .QN());
   DFF_X1 \MEM_reg[14][4]  (.D(n_32_20), .CK(n_32_1), .Q(\MEM[14] [4]), .QN());
   DFF_X1 \MEM_reg[14][3]  (.D(n_32_19), .CK(n_32_1), .Q(\MEM[14] [3]), .QN());
   DFF_X1 \MEM_reg[14][2]  (.D(n_32_18), .CK(n_32_1), .Q(\MEM[14] [2]), .QN());
   DFF_X1 \MEM_reg[14][1]  (.D(n_32_17), .CK(n_32_1), .Q(\MEM[14] [1]), .QN());
   DFF_X1 \MEM_reg[14][0]  (.D(n_32_16), .CK(n_32_1), .Q(\MEM[14] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[13]_reg  (.CK(clk), .E(n_32_61), .SE(1'b0), 
      .GCK(n_32_2));
   DFF_X1 \MEM_reg[13][31]  (.D(n_32_47), .CK(n_32_2), .Q(\MEM[13] [31]), .QN());
   DFF_X1 \MEM_reg[13][30]  (.D(n_32_46), .CK(n_32_2), .Q(\MEM[13] [30]), .QN());
   DFF_X1 \MEM_reg[13][29]  (.D(n_32_45), .CK(n_32_2), .Q(\MEM[13] [29]), .QN());
   DFF_X1 \MEM_reg[13][28]  (.D(n_32_44), .CK(n_32_2), .Q(\MEM[13] [28]), .QN());
   DFF_X1 \MEM_reg[13][27]  (.D(n_32_43), .CK(n_32_2), .Q(\MEM[13] [27]), .QN());
   DFF_X1 \MEM_reg[13][26]  (.D(n_32_42), .CK(n_32_2), .Q(\MEM[13] [26]), .QN());
   DFF_X1 \MEM_reg[13][25]  (.D(n_32_41), .CK(n_32_2), .Q(\MEM[13] [25]), .QN());
   DFF_X1 \MEM_reg[13][24]  (.D(n_32_40), .CK(n_32_2), .Q(\MEM[13] [24]), .QN());
   DFF_X1 \MEM_reg[13][23]  (.D(n_32_39), .CK(n_32_2), .Q(\MEM[13] [23]), .QN());
   DFF_X1 \MEM_reg[13][22]  (.D(n_32_38), .CK(n_32_2), .Q(\MEM[13] [22]), .QN());
   DFF_X1 \MEM_reg[13][21]  (.D(n_32_37), .CK(n_32_2), .Q(\MEM[13] [21]), .QN());
   DFF_X1 \MEM_reg[13][20]  (.D(n_32_36), .CK(n_32_2), .Q(\MEM[13] [20]), .QN());
   DFF_X1 \MEM_reg[13][19]  (.D(n_32_35), .CK(n_32_2), .Q(\MEM[13] [19]), .QN());
   DFF_X1 \MEM_reg[13][18]  (.D(n_32_34), .CK(n_32_2), .Q(\MEM[13] [18]), .QN());
   DFF_X1 \MEM_reg[13][17]  (.D(n_32_33), .CK(n_32_2), .Q(\MEM[13] [17]), .QN());
   DFF_X1 \MEM_reg[13][16]  (.D(n_32_32), .CK(n_32_2), .Q(\MEM[13] [16]), .QN());
   DFF_X1 \MEM_reg[13][15]  (.D(n_32_31), .CK(n_32_2), .Q(\MEM[13] [15]), .QN());
   DFF_X1 \MEM_reg[13][14]  (.D(n_32_30), .CK(n_32_2), .Q(\MEM[13] [14]), .QN());
   DFF_X1 \MEM_reg[13][13]  (.D(n_32_29), .CK(n_32_2), .Q(\MEM[13] [13]), .QN());
   DFF_X1 \MEM_reg[13][12]  (.D(n_32_28), .CK(n_32_2), .Q(\MEM[13] [12]), .QN());
   DFF_X1 \MEM_reg[13][11]  (.D(n_32_27), .CK(n_32_2), .Q(\MEM[13] [11]), .QN());
   DFF_X1 \MEM_reg[13][10]  (.D(n_32_26), .CK(n_32_2), .Q(\MEM[13] [10]), .QN());
   DFF_X1 \MEM_reg[13][9]  (.D(n_32_25), .CK(n_32_2), .Q(\MEM[13] [9]), .QN());
   DFF_X1 \MEM_reg[13][8]  (.D(n_32_24), .CK(n_32_2), .Q(\MEM[13] [8]), .QN());
   DFF_X1 \MEM_reg[13][7]  (.D(n_32_23), .CK(n_32_2), .Q(\MEM[13] [7]), .QN());
   DFF_X1 \MEM_reg[13][6]  (.D(n_32_22), .CK(n_32_2), .Q(\MEM[13] [6]), .QN());
   DFF_X1 \MEM_reg[13][5]  (.D(n_32_21), .CK(n_32_2), .Q(\MEM[13] [5]), .QN());
   DFF_X1 \MEM_reg[13][4]  (.D(n_32_20), .CK(n_32_2), .Q(\MEM[13] [4]), .QN());
   DFF_X1 \MEM_reg[13][3]  (.D(n_32_19), .CK(n_32_2), .Q(\MEM[13] [3]), .QN());
   DFF_X1 \MEM_reg[13][2]  (.D(n_32_18), .CK(n_32_2), .Q(\MEM[13] [2]), .QN());
   DFF_X1 \MEM_reg[13][1]  (.D(n_32_17), .CK(n_32_2), .Q(\MEM[13] [1]), .QN());
   DFF_X1 \MEM_reg[13][0]  (.D(n_32_16), .CK(n_32_2), .Q(\MEM[13] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[12]_reg  (.CK(clk), .E(n_32_60), .SE(1'b0), 
      .GCK(n_32_3));
   DFF_X1 \MEM_reg[12][31]  (.D(n_32_47), .CK(n_32_3), .Q(\MEM[12] [31]), .QN());
   DFF_X1 \MEM_reg[12][30]  (.D(n_32_46), .CK(n_32_3), .Q(\MEM[12] [30]), .QN());
   DFF_X1 \MEM_reg[12][29]  (.D(n_32_45), .CK(n_32_3), .Q(\MEM[12] [29]), .QN());
   DFF_X1 \MEM_reg[12][28]  (.D(n_32_44), .CK(n_32_3), .Q(\MEM[12] [28]), .QN());
   DFF_X1 \MEM_reg[12][27]  (.D(n_32_43), .CK(n_32_3), .Q(\MEM[12] [27]), .QN());
   DFF_X1 \MEM_reg[12][26]  (.D(n_32_42), .CK(n_32_3), .Q(\MEM[12] [26]), .QN());
   DFF_X1 \MEM_reg[12][25]  (.D(n_32_41), .CK(n_32_3), .Q(\MEM[12] [25]), .QN());
   DFF_X1 \MEM_reg[12][24]  (.D(n_32_40), .CK(n_32_3), .Q(\MEM[12] [24]), .QN());
   DFF_X1 \MEM_reg[12][23]  (.D(n_32_39), .CK(n_32_3), .Q(\MEM[12] [23]), .QN());
   DFF_X1 \MEM_reg[12][22]  (.D(n_32_38), .CK(n_32_3), .Q(\MEM[12] [22]), .QN());
   DFF_X1 \MEM_reg[12][21]  (.D(n_32_37), .CK(n_32_3), .Q(\MEM[12] [21]), .QN());
   DFF_X1 \MEM_reg[12][20]  (.D(n_32_36), .CK(n_32_3), .Q(\MEM[12] [20]), .QN());
   DFF_X1 \MEM_reg[12][19]  (.D(n_32_35), .CK(n_32_3), .Q(\MEM[12] [19]), .QN());
   DFF_X1 \MEM_reg[12][18]  (.D(n_32_34), .CK(n_32_3), .Q(\MEM[12] [18]), .QN());
   DFF_X1 \MEM_reg[12][17]  (.D(n_32_33), .CK(n_32_3), .Q(\MEM[12] [17]), .QN());
   DFF_X1 \MEM_reg[12][16]  (.D(n_32_32), .CK(n_32_3), .Q(\MEM[12] [16]), .QN());
   DFF_X1 \MEM_reg[12][15]  (.D(n_32_31), .CK(n_32_3), .Q(\MEM[12] [15]), .QN());
   DFF_X1 \MEM_reg[12][14]  (.D(n_32_30), .CK(n_32_3), .Q(\MEM[12] [14]), .QN());
   DFF_X1 \MEM_reg[12][13]  (.D(n_32_29), .CK(n_32_3), .Q(\MEM[12] [13]), .QN());
   DFF_X1 \MEM_reg[12][12]  (.D(n_32_28), .CK(n_32_3), .Q(\MEM[12] [12]), .QN());
   DFF_X1 \MEM_reg[12][11]  (.D(n_32_27), .CK(n_32_3), .Q(\MEM[12] [11]), .QN());
   DFF_X1 \MEM_reg[12][10]  (.D(n_32_26), .CK(n_32_3), .Q(\MEM[12] [10]), .QN());
   DFF_X1 \MEM_reg[12][9]  (.D(n_32_25), .CK(n_32_3), .Q(\MEM[12] [9]), .QN());
   DFF_X1 \MEM_reg[12][8]  (.D(n_32_24), .CK(n_32_3), .Q(\MEM[12] [8]), .QN());
   DFF_X1 \MEM_reg[12][7]  (.D(n_32_23), .CK(n_32_3), .Q(\MEM[12] [7]), .QN());
   DFF_X1 \MEM_reg[12][6]  (.D(n_32_22), .CK(n_32_3), .Q(\MEM[12] [6]), .QN());
   DFF_X1 \MEM_reg[12][5]  (.D(n_32_21), .CK(n_32_3), .Q(\MEM[12] [5]), .QN());
   DFF_X1 \MEM_reg[12][4]  (.D(n_32_20), .CK(n_32_3), .Q(\MEM[12] [4]), .QN());
   DFF_X1 \MEM_reg[12][3]  (.D(n_32_19), .CK(n_32_3), .Q(\MEM[12] [3]), .QN());
   DFF_X1 \MEM_reg[12][2]  (.D(n_32_18), .CK(n_32_3), .Q(\MEM[12] [2]), .QN());
   DFF_X1 \MEM_reg[12][1]  (.D(n_32_17), .CK(n_32_3), .Q(\MEM[12] [1]), .QN());
   DFF_X1 \MEM_reg[12][0]  (.D(n_32_16), .CK(n_32_3), .Q(\MEM[12] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[11]_reg  (.CK(clk), .E(n_32_59), .SE(1'b0), 
      .GCK(n_32_4));
   DFF_X1 \MEM_reg[11][31]  (.D(n_32_47), .CK(n_32_4), .Q(\MEM[11] [31]), .QN());
   DFF_X1 \MEM_reg[11][30]  (.D(n_32_46), .CK(n_32_4), .Q(\MEM[11] [30]), .QN());
   DFF_X1 \MEM_reg[11][29]  (.D(n_32_45), .CK(n_32_4), .Q(\MEM[11] [29]), .QN());
   DFF_X1 \MEM_reg[11][28]  (.D(n_32_44), .CK(n_32_4), .Q(\MEM[11] [28]), .QN());
   DFF_X1 \MEM_reg[11][27]  (.D(n_32_43), .CK(n_32_4), .Q(\MEM[11] [27]), .QN());
   DFF_X1 \MEM_reg[11][26]  (.D(n_32_42), .CK(n_32_4), .Q(\MEM[11] [26]), .QN());
   DFF_X1 \MEM_reg[11][25]  (.D(n_32_41), .CK(n_32_4), .Q(\MEM[11] [25]), .QN());
   DFF_X1 \MEM_reg[11][24]  (.D(n_32_40), .CK(n_32_4), .Q(\MEM[11] [24]), .QN());
   DFF_X1 \MEM_reg[11][23]  (.D(n_32_39), .CK(n_32_4), .Q(\MEM[11] [23]), .QN());
   DFF_X1 \MEM_reg[11][22]  (.D(n_32_38), .CK(n_32_4), .Q(\MEM[11] [22]), .QN());
   DFF_X1 \MEM_reg[11][21]  (.D(n_32_37), .CK(n_32_4), .Q(\MEM[11] [21]), .QN());
   DFF_X1 \MEM_reg[11][20]  (.D(n_32_36), .CK(n_32_4), .Q(\MEM[11] [20]), .QN());
   DFF_X1 \MEM_reg[11][19]  (.D(n_32_35), .CK(n_32_4), .Q(\MEM[11] [19]), .QN());
   DFF_X1 \MEM_reg[11][18]  (.D(n_32_34), .CK(n_32_4), .Q(\MEM[11] [18]), .QN());
   DFF_X1 \MEM_reg[11][17]  (.D(n_32_33), .CK(n_32_4), .Q(\MEM[11] [17]), .QN());
   DFF_X1 \MEM_reg[11][16]  (.D(n_32_32), .CK(n_32_4), .Q(\MEM[11] [16]), .QN());
   DFF_X1 \MEM_reg[11][15]  (.D(n_32_31), .CK(n_32_4), .Q(\MEM[11] [15]), .QN());
   DFF_X1 \MEM_reg[11][14]  (.D(n_32_30), .CK(n_32_4), .Q(\MEM[11] [14]), .QN());
   DFF_X1 \MEM_reg[11][13]  (.D(n_32_29), .CK(n_32_4), .Q(\MEM[11] [13]), .QN());
   DFF_X1 \MEM_reg[11][12]  (.D(n_32_28), .CK(n_32_4), .Q(\MEM[11] [12]), .QN());
   DFF_X1 \MEM_reg[11][11]  (.D(n_32_27), .CK(n_32_4), .Q(\MEM[11] [11]), .QN());
   DFF_X1 \MEM_reg[11][10]  (.D(n_32_26), .CK(n_32_4), .Q(\MEM[11] [10]), .QN());
   DFF_X1 \MEM_reg[11][9]  (.D(n_32_25), .CK(n_32_4), .Q(\MEM[11] [9]), .QN());
   DFF_X1 \MEM_reg[11][8]  (.D(n_32_24), .CK(n_32_4), .Q(\MEM[11] [8]), .QN());
   DFF_X1 \MEM_reg[11][7]  (.D(n_32_23), .CK(n_32_4), .Q(\MEM[11] [7]), .QN());
   DFF_X1 \MEM_reg[11][6]  (.D(n_32_22), .CK(n_32_4), .Q(\MEM[11] [6]), .QN());
   DFF_X1 \MEM_reg[11][5]  (.D(n_32_21), .CK(n_32_4), .Q(\MEM[11] [5]), .QN());
   DFF_X1 \MEM_reg[11][4]  (.D(n_32_20), .CK(n_32_4), .Q(\MEM[11] [4]), .QN());
   DFF_X1 \MEM_reg[11][3]  (.D(n_32_19), .CK(n_32_4), .Q(\MEM[11] [3]), .QN());
   DFF_X1 \MEM_reg[11][2]  (.D(n_32_18), .CK(n_32_4), .Q(\MEM[11] [2]), .QN());
   DFF_X1 \MEM_reg[11][1]  (.D(n_32_17), .CK(n_32_4), .Q(\MEM[11] [1]), .QN());
   DFF_X1 \MEM_reg[11][0]  (.D(n_32_16), .CK(n_32_4), .Q(\MEM[11] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[10]_reg  (.CK(clk), .E(n_32_58), .SE(1'b0), 
      .GCK(n_32_5));
   DFF_X1 \MEM_reg[10][31]  (.D(n_32_47), .CK(n_32_5), .Q(\MEM[10] [31]), .QN());
   DFF_X1 \MEM_reg[10][30]  (.D(n_32_46), .CK(n_32_5), .Q(\MEM[10] [30]), .QN());
   DFF_X1 \MEM_reg[10][29]  (.D(n_32_45), .CK(n_32_5), .Q(\MEM[10] [29]), .QN());
   DFF_X1 \MEM_reg[10][28]  (.D(n_32_44), .CK(n_32_5), .Q(\MEM[10] [28]), .QN());
   DFF_X1 \MEM_reg[10][27]  (.D(n_32_43), .CK(n_32_5), .Q(\MEM[10] [27]), .QN());
   DFF_X1 \MEM_reg[10][26]  (.D(n_32_42), .CK(n_32_5), .Q(\MEM[10] [26]), .QN());
   DFF_X1 \MEM_reg[10][25]  (.D(n_32_41), .CK(n_32_5), .Q(\MEM[10] [25]), .QN());
   DFF_X1 \MEM_reg[10][24]  (.D(n_32_40), .CK(n_32_5), .Q(\MEM[10] [24]), .QN());
   DFF_X1 \MEM_reg[10][23]  (.D(n_32_39), .CK(n_32_5), .Q(\MEM[10] [23]), .QN());
   DFF_X1 \MEM_reg[10][22]  (.D(n_32_38), .CK(n_32_5), .Q(\MEM[10] [22]), .QN());
   DFF_X1 \MEM_reg[10][21]  (.D(n_32_37), .CK(n_32_5), .Q(\MEM[10] [21]), .QN());
   DFF_X1 \MEM_reg[10][20]  (.D(n_32_36), .CK(n_32_5), .Q(\MEM[10] [20]), .QN());
   DFF_X1 \MEM_reg[10][19]  (.D(n_32_35), .CK(n_32_5), .Q(\MEM[10] [19]), .QN());
   DFF_X1 \MEM_reg[10][18]  (.D(n_32_34), .CK(n_32_5), .Q(\MEM[10] [18]), .QN());
   DFF_X1 \MEM_reg[10][17]  (.D(n_32_33), .CK(n_32_5), .Q(\MEM[10] [17]), .QN());
   DFF_X1 \MEM_reg[10][16]  (.D(n_32_32), .CK(n_32_5), .Q(\MEM[10] [16]), .QN());
   DFF_X1 \MEM_reg[10][15]  (.D(n_32_31), .CK(n_32_5), .Q(\MEM[10] [15]), .QN());
   DFF_X1 \MEM_reg[10][14]  (.D(n_32_30), .CK(n_32_5), .Q(\MEM[10] [14]), .QN());
   DFF_X1 \MEM_reg[10][13]  (.D(n_32_29), .CK(n_32_5), .Q(\MEM[10] [13]), .QN());
   DFF_X1 \MEM_reg[10][12]  (.D(n_32_28), .CK(n_32_5), .Q(\MEM[10] [12]), .QN());
   DFF_X1 \MEM_reg[10][11]  (.D(n_32_27), .CK(n_32_5), .Q(\MEM[10] [11]), .QN());
   DFF_X1 \MEM_reg[10][10]  (.D(n_32_26), .CK(n_32_5), .Q(\MEM[10] [10]), .QN());
   DFF_X1 \MEM_reg[10][9]  (.D(n_32_25), .CK(n_32_5), .Q(\MEM[10] [9]), .QN());
   DFF_X1 \MEM_reg[10][8]  (.D(n_32_24), .CK(n_32_5), .Q(\MEM[10] [8]), .QN());
   DFF_X1 \MEM_reg[10][7]  (.D(n_32_23), .CK(n_32_5), .Q(\MEM[10] [7]), .QN());
   DFF_X1 \MEM_reg[10][6]  (.D(n_32_22), .CK(n_32_5), .Q(\MEM[10] [6]), .QN());
   DFF_X1 \MEM_reg[10][5]  (.D(n_32_21), .CK(n_32_5), .Q(\MEM[10] [5]), .QN());
   DFF_X1 \MEM_reg[10][4]  (.D(n_32_20), .CK(n_32_5), .Q(\MEM[10] [4]), .QN());
   DFF_X1 \MEM_reg[10][3]  (.D(n_32_19), .CK(n_32_5), .Q(\MEM[10] [3]), .QN());
   DFF_X1 \MEM_reg[10][2]  (.D(n_32_18), .CK(n_32_5), .Q(\MEM[10] [2]), .QN());
   DFF_X1 \MEM_reg[10][1]  (.D(n_32_17), .CK(n_32_5), .Q(\MEM[10] [1]), .QN());
   DFF_X1 \MEM_reg[10][0]  (.D(n_32_16), .CK(n_32_5), .Q(\MEM[10] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[9]_reg  (.CK(clk), .E(n_32_57), .SE(1'b0), 
      .GCK(n_32_6));
   DFF_X1 \MEM_reg[9][31]  (.D(n_32_47), .CK(n_32_6), .Q(\MEM[9] [31]), .QN());
   DFF_X1 \MEM_reg[9][30]  (.D(n_32_46), .CK(n_32_6), .Q(\MEM[9] [30]), .QN());
   DFF_X1 \MEM_reg[9][29]  (.D(n_32_45), .CK(n_32_6), .Q(\MEM[9] [29]), .QN());
   DFF_X1 \MEM_reg[9][28]  (.D(n_32_44), .CK(n_32_6), .Q(\MEM[9] [28]), .QN());
   DFF_X1 \MEM_reg[9][27]  (.D(n_32_43), .CK(n_32_6), .Q(\MEM[9] [27]), .QN());
   DFF_X1 \MEM_reg[9][26]  (.D(n_32_42), .CK(n_32_6), .Q(\MEM[9] [26]), .QN());
   DFF_X1 \MEM_reg[9][25]  (.D(n_32_41), .CK(n_32_6), .Q(\MEM[9] [25]), .QN());
   DFF_X1 \MEM_reg[9][24]  (.D(n_32_40), .CK(n_32_6), .Q(\MEM[9] [24]), .QN());
   DFF_X1 \MEM_reg[9][23]  (.D(n_32_39), .CK(n_32_6), .Q(\MEM[9] [23]), .QN());
   DFF_X1 \MEM_reg[9][22]  (.D(n_32_38), .CK(n_32_6), .Q(\MEM[9] [22]), .QN());
   DFF_X1 \MEM_reg[9][21]  (.D(n_32_37), .CK(n_32_6), .Q(\MEM[9] [21]), .QN());
   DFF_X1 \MEM_reg[9][20]  (.D(n_32_36), .CK(n_32_6), .Q(\MEM[9] [20]), .QN());
   DFF_X1 \MEM_reg[9][19]  (.D(n_32_35), .CK(n_32_6), .Q(\MEM[9] [19]), .QN());
   DFF_X1 \MEM_reg[9][18]  (.D(n_32_34), .CK(n_32_6), .Q(\MEM[9] [18]), .QN());
   DFF_X1 \MEM_reg[9][17]  (.D(n_32_33), .CK(n_32_6), .Q(\MEM[9] [17]), .QN());
   DFF_X1 \MEM_reg[9][16]  (.D(n_32_32), .CK(n_32_6), .Q(\MEM[9] [16]), .QN());
   DFF_X1 \MEM_reg[9][15]  (.D(n_32_31), .CK(n_32_6), .Q(\MEM[9] [15]), .QN());
   DFF_X1 \MEM_reg[9][14]  (.D(n_32_30), .CK(n_32_6), .Q(\MEM[9] [14]), .QN());
   DFF_X1 \MEM_reg[9][13]  (.D(n_32_29), .CK(n_32_6), .Q(\MEM[9] [13]), .QN());
   DFF_X1 \MEM_reg[9][12]  (.D(n_32_28), .CK(n_32_6), .Q(\MEM[9] [12]), .QN());
   DFF_X1 \MEM_reg[9][11]  (.D(n_32_27), .CK(n_32_6), .Q(\MEM[9] [11]), .QN());
   DFF_X1 \MEM_reg[9][10]  (.D(n_32_26), .CK(n_32_6), .Q(\MEM[9] [10]), .QN());
   DFF_X1 \MEM_reg[9][9]  (.D(n_32_25), .CK(n_32_6), .Q(\MEM[9] [9]), .QN());
   DFF_X1 \MEM_reg[9][8]  (.D(n_32_24), .CK(n_32_6), .Q(\MEM[9] [8]), .QN());
   DFF_X1 \MEM_reg[9][7]  (.D(n_32_23), .CK(n_32_6), .Q(\MEM[9] [7]), .QN());
   DFF_X1 \MEM_reg[9][6]  (.D(n_32_22), .CK(n_32_6), .Q(\MEM[9] [6]), .QN());
   DFF_X1 \MEM_reg[9][5]  (.D(n_32_21), .CK(n_32_6), .Q(\MEM[9] [5]), .QN());
   DFF_X1 \MEM_reg[9][4]  (.D(n_32_20), .CK(n_32_6), .Q(\MEM[9] [4]), .QN());
   DFF_X1 \MEM_reg[9][3]  (.D(n_32_19), .CK(n_32_6), .Q(\MEM[9] [3]), .QN());
   DFF_X1 \MEM_reg[9][2]  (.D(n_32_18), .CK(n_32_6), .Q(\MEM[9] [2]), .QN());
   DFF_X1 \MEM_reg[9][1]  (.D(n_32_17), .CK(n_32_6), .Q(\MEM[9] [1]), .QN());
   DFF_X1 \MEM_reg[9][0]  (.D(n_32_16), .CK(n_32_6), .Q(\MEM[9] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[8]_reg  (.CK(clk), .E(n_32_56), .SE(1'b0), 
      .GCK(n_32_7));
   DFF_X1 \MEM_reg[8][31]  (.D(n_32_47), .CK(n_32_7), .Q(\MEM[8] [31]), .QN());
   DFF_X1 \MEM_reg[8][30]  (.D(n_32_46), .CK(n_32_7), .Q(\MEM[8] [30]), .QN());
   DFF_X1 \MEM_reg[8][29]  (.D(n_32_45), .CK(n_32_7), .Q(\MEM[8] [29]), .QN());
   DFF_X1 \MEM_reg[8][28]  (.D(n_32_44), .CK(n_32_7), .Q(\MEM[8] [28]), .QN());
   DFF_X1 \MEM_reg[8][27]  (.D(n_32_43), .CK(n_32_7), .Q(\MEM[8] [27]), .QN());
   DFF_X1 \MEM_reg[8][26]  (.D(n_32_42), .CK(n_32_7), .Q(\MEM[8] [26]), .QN());
   DFF_X1 \MEM_reg[8][25]  (.D(n_32_41), .CK(n_32_7), .Q(\MEM[8] [25]), .QN());
   DFF_X1 \MEM_reg[8][24]  (.D(n_32_40), .CK(n_32_7), .Q(\MEM[8] [24]), .QN());
   DFF_X1 \MEM_reg[8][23]  (.D(n_32_39), .CK(n_32_7), .Q(\MEM[8] [23]), .QN());
   DFF_X1 \MEM_reg[8][22]  (.D(n_32_38), .CK(n_32_7), .Q(\MEM[8] [22]), .QN());
   DFF_X1 \MEM_reg[8][21]  (.D(n_32_37), .CK(n_32_7), .Q(\MEM[8] [21]), .QN());
   DFF_X1 \MEM_reg[8][20]  (.D(n_32_36), .CK(n_32_7), .Q(\MEM[8] [20]), .QN());
   DFF_X1 \MEM_reg[8][19]  (.D(n_32_35), .CK(n_32_7), .Q(\MEM[8] [19]), .QN());
   DFF_X1 \MEM_reg[8][18]  (.D(n_32_34), .CK(n_32_7), .Q(\MEM[8] [18]), .QN());
   DFF_X1 \MEM_reg[8][17]  (.D(n_32_33), .CK(n_32_7), .Q(\MEM[8] [17]), .QN());
   DFF_X1 \MEM_reg[8][16]  (.D(n_32_32), .CK(n_32_7), .Q(\MEM[8] [16]), .QN());
   DFF_X1 \MEM_reg[8][15]  (.D(n_32_31), .CK(n_32_7), .Q(\MEM[8] [15]), .QN());
   DFF_X1 \MEM_reg[8][14]  (.D(n_32_30), .CK(n_32_7), .Q(\MEM[8] [14]), .QN());
   DFF_X1 \MEM_reg[8][13]  (.D(n_32_29), .CK(n_32_7), .Q(\MEM[8] [13]), .QN());
   DFF_X1 \MEM_reg[8][12]  (.D(n_32_28), .CK(n_32_7), .Q(\MEM[8] [12]), .QN());
   DFF_X1 \MEM_reg[8][11]  (.D(n_32_27), .CK(n_32_7), .Q(\MEM[8] [11]), .QN());
   DFF_X1 \MEM_reg[8][10]  (.D(n_32_26), .CK(n_32_7), .Q(\MEM[8] [10]), .QN());
   DFF_X1 \MEM_reg[8][9]  (.D(n_32_25), .CK(n_32_7), .Q(\MEM[8] [9]), .QN());
   DFF_X1 \MEM_reg[8][8]  (.D(n_32_24), .CK(n_32_7), .Q(\MEM[8] [8]), .QN());
   DFF_X1 \MEM_reg[8][7]  (.D(n_32_23), .CK(n_32_7), .Q(\MEM[8] [7]), .QN());
   DFF_X1 \MEM_reg[8][6]  (.D(n_32_22), .CK(n_32_7), .Q(\MEM[8] [6]), .QN());
   DFF_X1 \MEM_reg[8][5]  (.D(n_32_21), .CK(n_32_7), .Q(\MEM[8] [5]), .QN());
   DFF_X1 \MEM_reg[8][4]  (.D(n_32_20), .CK(n_32_7), .Q(\MEM[8] [4]), .QN());
   DFF_X1 \MEM_reg[8][3]  (.D(n_32_19), .CK(n_32_7), .Q(\MEM[8] [3]), .QN());
   DFF_X1 \MEM_reg[8][2]  (.D(n_32_18), .CK(n_32_7), .Q(\MEM[8] [2]), .QN());
   DFF_X1 \MEM_reg[8][1]  (.D(n_32_17), .CK(n_32_7), .Q(\MEM[8] [1]), .QN());
   DFF_X1 \MEM_reg[8][0]  (.D(n_32_16), .CK(n_32_7), .Q(\MEM[8] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[7]_reg  (.CK(clk), .E(n_32_55), .SE(1'b0), 
      .GCK(n_32_8));
   DFF_X1 \MEM_reg[7][31]  (.D(n_32_47), .CK(n_32_8), .Q(\MEM[7] [31]), .QN());
   DFF_X1 \MEM_reg[7][30]  (.D(n_32_46), .CK(n_32_8), .Q(\MEM[7] [30]), .QN());
   DFF_X1 \MEM_reg[7][29]  (.D(n_32_45), .CK(n_32_8), .Q(\MEM[7] [29]), .QN());
   DFF_X1 \MEM_reg[7][28]  (.D(n_32_44), .CK(n_32_8), .Q(\MEM[7] [28]), .QN());
   DFF_X1 \MEM_reg[7][27]  (.D(n_32_43), .CK(n_32_8), .Q(\MEM[7] [27]), .QN());
   DFF_X1 \MEM_reg[7][26]  (.D(n_32_42), .CK(n_32_8), .Q(\MEM[7] [26]), .QN());
   DFF_X1 \MEM_reg[7][25]  (.D(n_32_41), .CK(n_32_8), .Q(\MEM[7] [25]), .QN());
   DFF_X1 \MEM_reg[7][24]  (.D(n_32_40), .CK(n_32_8), .Q(\MEM[7] [24]), .QN());
   DFF_X1 \MEM_reg[7][23]  (.D(n_32_39), .CK(n_32_8), .Q(\MEM[7] [23]), .QN());
   DFF_X1 \MEM_reg[7][22]  (.D(n_32_38), .CK(n_32_8), .Q(\MEM[7] [22]), .QN());
   DFF_X1 \MEM_reg[7][21]  (.D(n_32_37), .CK(n_32_8), .Q(\MEM[7] [21]), .QN());
   DFF_X1 \MEM_reg[7][20]  (.D(n_32_36), .CK(n_32_8), .Q(\MEM[7] [20]), .QN());
   DFF_X1 \MEM_reg[7][19]  (.D(n_32_35), .CK(n_32_8), .Q(\MEM[7] [19]), .QN());
   DFF_X1 \MEM_reg[7][18]  (.D(n_32_34), .CK(n_32_8), .Q(\MEM[7] [18]), .QN());
   DFF_X1 \MEM_reg[7][17]  (.D(n_32_33), .CK(n_32_8), .Q(\MEM[7] [17]), .QN());
   DFF_X1 \MEM_reg[7][16]  (.D(n_32_32), .CK(n_32_8), .Q(\MEM[7] [16]), .QN());
   DFF_X1 \MEM_reg[7][15]  (.D(n_32_31), .CK(n_32_8), .Q(\MEM[7] [15]), .QN());
   DFF_X1 \MEM_reg[7][14]  (.D(n_32_30), .CK(n_32_8), .Q(\MEM[7] [14]), .QN());
   DFF_X1 \MEM_reg[7][13]  (.D(n_32_29), .CK(n_32_8), .Q(\MEM[7] [13]), .QN());
   DFF_X1 \MEM_reg[7][12]  (.D(n_32_28), .CK(n_32_8), .Q(\MEM[7] [12]), .QN());
   DFF_X1 \MEM_reg[7][11]  (.D(n_32_27), .CK(n_32_8), .Q(\MEM[7] [11]), .QN());
   DFF_X1 \MEM_reg[7][10]  (.D(n_32_26), .CK(n_32_8), .Q(\MEM[7] [10]), .QN());
   DFF_X1 \MEM_reg[7][9]  (.D(n_32_25), .CK(n_32_8), .Q(\MEM[7] [9]), .QN());
   DFF_X1 \MEM_reg[7][8]  (.D(n_32_24), .CK(n_32_8), .Q(\MEM[7] [8]), .QN());
   DFF_X1 \MEM_reg[7][7]  (.D(n_32_23), .CK(n_32_8), .Q(\MEM[7] [7]), .QN());
   DFF_X1 \MEM_reg[7][6]  (.D(n_32_22), .CK(n_32_8), .Q(\MEM[7] [6]), .QN());
   DFF_X1 \MEM_reg[7][5]  (.D(n_32_21), .CK(n_32_8), .Q(\MEM[7] [5]), .QN());
   DFF_X1 \MEM_reg[7][4]  (.D(n_32_20), .CK(n_32_8), .Q(\MEM[7] [4]), .QN());
   DFF_X1 \MEM_reg[7][3]  (.D(n_32_19), .CK(n_32_8), .Q(\MEM[7] [3]), .QN());
   DFF_X1 \MEM_reg[7][2]  (.D(n_32_18), .CK(n_32_8), .Q(\MEM[7] [2]), .QN());
   DFF_X1 \MEM_reg[7][1]  (.D(n_32_17), .CK(n_32_8), .Q(\MEM[7] [1]), .QN());
   DFF_X1 \MEM_reg[7][0]  (.D(n_32_16), .CK(n_32_8), .Q(\MEM[7] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[6]_reg  (.CK(clk), .E(n_32_54), .SE(1'b0), 
      .GCK(n_32_9));
   DFF_X1 \MEM_reg[6][31]  (.D(n_32_47), .CK(n_32_9), .Q(\MEM[6] [31]), .QN());
   DFF_X1 \MEM_reg[6][30]  (.D(n_32_46), .CK(n_32_9), .Q(\MEM[6] [30]), .QN());
   DFF_X1 \MEM_reg[6][29]  (.D(n_32_45), .CK(n_32_9), .Q(\MEM[6] [29]), .QN());
   DFF_X1 \MEM_reg[6][28]  (.D(n_32_44), .CK(n_32_9), .Q(\MEM[6] [28]), .QN());
   DFF_X1 \MEM_reg[6][27]  (.D(n_32_43), .CK(n_32_9), .Q(\MEM[6] [27]), .QN());
   DFF_X1 \MEM_reg[6][26]  (.D(n_32_42), .CK(n_32_9), .Q(\MEM[6] [26]), .QN());
   DFF_X1 \MEM_reg[6][25]  (.D(n_32_41), .CK(n_32_9), .Q(\MEM[6] [25]), .QN());
   DFF_X1 \MEM_reg[6][24]  (.D(n_32_40), .CK(n_32_9), .Q(\MEM[6] [24]), .QN());
   DFF_X1 \MEM_reg[6][23]  (.D(n_32_39), .CK(n_32_9), .Q(\MEM[6] [23]), .QN());
   DFF_X1 \MEM_reg[6][22]  (.D(n_32_38), .CK(n_32_9), .Q(\MEM[6] [22]), .QN());
   DFF_X1 \MEM_reg[6][21]  (.D(n_32_37), .CK(n_32_9), .Q(\MEM[6] [21]), .QN());
   DFF_X1 \MEM_reg[6][20]  (.D(n_32_36), .CK(n_32_9), .Q(\MEM[6] [20]), .QN());
   DFF_X1 \MEM_reg[6][19]  (.D(n_32_35), .CK(n_32_9), .Q(\MEM[6] [19]), .QN());
   DFF_X1 \MEM_reg[6][18]  (.D(n_32_34), .CK(n_32_9), .Q(\MEM[6] [18]), .QN());
   DFF_X1 \MEM_reg[6][17]  (.D(n_32_33), .CK(n_32_9), .Q(\MEM[6] [17]), .QN());
   DFF_X1 \MEM_reg[6][16]  (.D(n_32_32), .CK(n_32_9), .Q(\MEM[6] [16]), .QN());
   DFF_X1 \MEM_reg[6][15]  (.D(n_32_31), .CK(n_32_9), .Q(\MEM[6] [15]), .QN());
   DFF_X1 \MEM_reg[6][14]  (.D(n_32_30), .CK(n_32_9), .Q(\MEM[6] [14]), .QN());
   DFF_X1 \MEM_reg[6][13]  (.D(n_32_29), .CK(n_32_9), .Q(\MEM[6] [13]), .QN());
   DFF_X1 \MEM_reg[6][12]  (.D(n_32_28), .CK(n_32_9), .Q(\MEM[6] [12]), .QN());
   DFF_X1 \MEM_reg[6][11]  (.D(n_32_27), .CK(n_32_9), .Q(\MEM[6] [11]), .QN());
   DFF_X1 \MEM_reg[6][10]  (.D(n_32_26), .CK(n_32_9), .Q(\MEM[6] [10]), .QN());
   DFF_X1 \MEM_reg[6][9]  (.D(n_32_25), .CK(n_32_9), .Q(\MEM[6] [9]), .QN());
   DFF_X1 \MEM_reg[6][8]  (.D(n_32_24), .CK(n_32_9), .Q(\MEM[6] [8]), .QN());
   DFF_X1 \MEM_reg[6][7]  (.D(n_32_23), .CK(n_32_9), .Q(\MEM[6] [7]), .QN());
   DFF_X1 \MEM_reg[6][6]  (.D(n_32_22), .CK(n_32_9), .Q(\MEM[6] [6]), .QN());
   DFF_X1 \MEM_reg[6][5]  (.D(n_32_21), .CK(n_32_9), .Q(\MEM[6] [5]), .QN());
   DFF_X1 \MEM_reg[6][4]  (.D(n_32_20), .CK(n_32_9), .Q(\MEM[6] [4]), .QN());
   DFF_X1 \MEM_reg[6][3]  (.D(n_32_19), .CK(n_32_9), .Q(\MEM[6] [3]), .QN());
   DFF_X1 \MEM_reg[6][2]  (.D(n_32_18), .CK(n_32_9), .Q(\MEM[6] [2]), .QN());
   DFF_X1 \MEM_reg[6][1]  (.D(n_32_17), .CK(n_32_9), .Q(\MEM[6] [1]), .QN());
   DFF_X1 \MEM_reg[6][0]  (.D(n_32_16), .CK(n_32_9), .Q(\MEM[6] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[5]_reg  (.CK(clk), .E(n_32_53), .SE(1'b0), 
      .GCK(n_32_10));
   DFF_X1 \MEM_reg[5][31]  (.D(n_32_47), .CK(n_32_10), .Q(\MEM[5] [31]), .QN());
   DFF_X1 \MEM_reg[5][30]  (.D(n_32_46), .CK(n_32_10), .Q(\MEM[5] [30]), .QN());
   DFF_X1 \MEM_reg[5][29]  (.D(n_32_45), .CK(n_32_10), .Q(\MEM[5] [29]), .QN());
   DFF_X1 \MEM_reg[5][28]  (.D(n_32_44), .CK(n_32_10), .Q(\MEM[5] [28]), .QN());
   DFF_X1 \MEM_reg[5][27]  (.D(n_32_43), .CK(n_32_10), .Q(\MEM[5] [27]), .QN());
   DFF_X1 \MEM_reg[5][26]  (.D(n_32_42), .CK(n_32_10), .Q(\MEM[5] [26]), .QN());
   DFF_X1 \MEM_reg[5][25]  (.D(n_32_41), .CK(n_32_10), .Q(\MEM[5] [25]), .QN());
   DFF_X1 \MEM_reg[5][24]  (.D(n_32_40), .CK(n_32_10), .Q(\MEM[5] [24]), .QN());
   DFF_X1 \MEM_reg[5][23]  (.D(n_32_39), .CK(n_32_10), .Q(\MEM[5] [23]), .QN());
   DFF_X1 \MEM_reg[5][22]  (.D(n_32_38), .CK(n_32_10), .Q(\MEM[5] [22]), .QN());
   DFF_X1 \MEM_reg[5][21]  (.D(n_32_37), .CK(n_32_10), .Q(\MEM[5] [21]), .QN());
   DFF_X1 \MEM_reg[5][20]  (.D(n_32_36), .CK(n_32_10), .Q(\MEM[5] [20]), .QN());
   DFF_X1 \MEM_reg[5][19]  (.D(n_32_35), .CK(n_32_10), .Q(\MEM[5] [19]), .QN());
   DFF_X1 \MEM_reg[5][18]  (.D(n_32_34), .CK(n_32_10), .Q(\MEM[5] [18]), .QN());
   DFF_X1 \MEM_reg[5][17]  (.D(n_32_33), .CK(n_32_10), .Q(\MEM[5] [17]), .QN());
   DFF_X1 \MEM_reg[5][16]  (.D(n_32_32), .CK(n_32_10), .Q(\MEM[5] [16]), .QN());
   DFF_X1 \MEM_reg[5][15]  (.D(n_32_31), .CK(n_32_10), .Q(\MEM[5] [15]), .QN());
   DFF_X1 \MEM_reg[5][14]  (.D(n_32_30), .CK(n_32_10), .Q(\MEM[5] [14]), .QN());
   DFF_X1 \MEM_reg[5][13]  (.D(n_32_29), .CK(n_32_10), .Q(\MEM[5] [13]), .QN());
   DFF_X1 \MEM_reg[5][12]  (.D(n_32_28), .CK(n_32_10), .Q(\MEM[5] [12]), .QN());
   DFF_X1 \MEM_reg[5][11]  (.D(n_32_27), .CK(n_32_10), .Q(\MEM[5] [11]), .QN());
   DFF_X1 \MEM_reg[5][10]  (.D(n_32_26), .CK(n_32_10), .Q(\MEM[5] [10]), .QN());
   DFF_X1 \MEM_reg[5][9]  (.D(n_32_25), .CK(n_32_10), .Q(\MEM[5] [9]), .QN());
   DFF_X1 \MEM_reg[5][8]  (.D(n_32_24), .CK(n_32_10), .Q(\MEM[5] [8]), .QN());
   DFF_X1 \MEM_reg[5][7]  (.D(n_32_23), .CK(n_32_10), .Q(\MEM[5] [7]), .QN());
   DFF_X1 \MEM_reg[5][6]  (.D(n_32_22), .CK(n_32_10), .Q(\MEM[5] [6]), .QN());
   DFF_X1 \MEM_reg[5][5]  (.D(n_32_21), .CK(n_32_10), .Q(\MEM[5] [5]), .QN());
   DFF_X1 \MEM_reg[5][4]  (.D(n_32_20), .CK(n_32_10), .Q(\MEM[5] [4]), .QN());
   DFF_X1 \MEM_reg[5][3]  (.D(n_32_19), .CK(n_32_10), .Q(\MEM[5] [3]), .QN());
   DFF_X1 \MEM_reg[5][2]  (.D(n_32_18), .CK(n_32_10), .Q(\MEM[5] [2]), .QN());
   DFF_X1 \MEM_reg[5][1]  (.D(n_32_17), .CK(n_32_10), .Q(\MEM[5] [1]), .QN());
   DFF_X1 \MEM_reg[5][0]  (.D(n_32_16), .CK(n_32_10), .Q(\MEM[5] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[4]_reg  (.CK(clk), .E(n_32_52), .SE(1'b0), 
      .GCK(n_32_11));
   DFF_X1 \MEM_reg[4][31]  (.D(n_32_47), .CK(n_32_11), .Q(\MEM[4] [31]), .QN());
   DFF_X1 \MEM_reg[4][30]  (.D(n_32_46), .CK(n_32_11), .Q(\MEM[4] [30]), .QN());
   DFF_X1 \MEM_reg[4][29]  (.D(n_32_45), .CK(n_32_11), .Q(\MEM[4] [29]), .QN());
   DFF_X1 \MEM_reg[4][28]  (.D(n_32_44), .CK(n_32_11), .Q(\MEM[4] [28]), .QN());
   DFF_X1 \MEM_reg[4][27]  (.D(n_32_43), .CK(n_32_11), .Q(\MEM[4] [27]), .QN());
   DFF_X1 \MEM_reg[4][26]  (.D(n_32_42), .CK(n_32_11), .Q(\MEM[4] [26]), .QN());
   DFF_X1 \MEM_reg[4][25]  (.D(n_32_41), .CK(n_32_11), .Q(\MEM[4] [25]), .QN());
   DFF_X1 \MEM_reg[4][24]  (.D(n_32_40), .CK(n_32_11), .Q(\MEM[4] [24]), .QN());
   DFF_X1 \MEM_reg[4][23]  (.D(n_32_39), .CK(n_32_11), .Q(\MEM[4] [23]), .QN());
   DFF_X1 \MEM_reg[4][22]  (.D(n_32_38), .CK(n_32_11), .Q(\MEM[4] [22]), .QN());
   DFF_X1 \MEM_reg[4][21]  (.D(n_32_37), .CK(n_32_11), .Q(\MEM[4] [21]), .QN());
   DFF_X1 \MEM_reg[4][20]  (.D(n_32_36), .CK(n_32_11), .Q(\MEM[4] [20]), .QN());
   DFF_X1 \MEM_reg[4][19]  (.D(n_32_35), .CK(n_32_11), .Q(\MEM[4] [19]), .QN());
   DFF_X1 \MEM_reg[4][18]  (.D(n_32_34), .CK(n_32_11), .Q(\MEM[4] [18]), .QN());
   DFF_X1 \MEM_reg[4][17]  (.D(n_32_33), .CK(n_32_11), .Q(\MEM[4] [17]), .QN());
   DFF_X1 \MEM_reg[4][16]  (.D(n_32_32), .CK(n_32_11), .Q(\MEM[4] [16]), .QN());
   DFF_X1 \MEM_reg[4][15]  (.D(n_32_31), .CK(n_32_11), .Q(\MEM[4] [15]), .QN());
   DFF_X1 \MEM_reg[4][14]  (.D(n_32_30), .CK(n_32_11), .Q(\MEM[4] [14]), .QN());
   DFF_X1 \MEM_reg[4][13]  (.D(n_32_29), .CK(n_32_11), .Q(\MEM[4] [13]), .QN());
   DFF_X1 \MEM_reg[4][12]  (.D(n_32_28), .CK(n_32_11), .Q(\MEM[4] [12]), .QN());
   DFF_X1 \MEM_reg[4][11]  (.D(n_32_27), .CK(n_32_11), .Q(\MEM[4] [11]), .QN());
   DFF_X1 \MEM_reg[4][10]  (.D(n_32_26), .CK(n_32_11), .Q(\MEM[4] [10]), .QN());
   DFF_X1 \MEM_reg[4][9]  (.D(n_32_25), .CK(n_32_11), .Q(\MEM[4] [9]), .QN());
   DFF_X1 \MEM_reg[4][8]  (.D(n_32_24), .CK(n_32_11), .Q(\MEM[4] [8]), .QN());
   DFF_X1 \MEM_reg[4][7]  (.D(n_32_23), .CK(n_32_11), .Q(\MEM[4] [7]), .QN());
   DFF_X1 \MEM_reg[4][6]  (.D(n_32_22), .CK(n_32_11), .Q(\MEM[4] [6]), .QN());
   DFF_X1 \MEM_reg[4][5]  (.D(n_32_21), .CK(n_32_11), .Q(\MEM[4] [5]), .QN());
   DFF_X1 \MEM_reg[4][4]  (.D(n_32_20), .CK(n_32_11), .Q(\MEM[4] [4]), .QN());
   DFF_X1 \MEM_reg[4][3]  (.D(n_32_19), .CK(n_32_11), .Q(\MEM[4] [3]), .QN());
   DFF_X1 \MEM_reg[4][2]  (.D(n_32_18), .CK(n_32_11), .Q(\MEM[4] [2]), .QN());
   DFF_X1 \MEM_reg[4][1]  (.D(n_32_17), .CK(n_32_11), .Q(\MEM[4] [1]), .QN());
   DFF_X1 \MEM_reg[4][0]  (.D(n_32_16), .CK(n_32_11), .Q(\MEM[4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[3]_reg  (.CK(clk), .E(n_32_51), .SE(1'b0), 
      .GCK(n_32_12));
   DFF_X1 \MEM_reg[3][31]  (.D(n_32_47), .CK(n_32_12), .Q(\MEM[3] [31]), .QN());
   DFF_X1 \MEM_reg[3][30]  (.D(n_32_46), .CK(n_32_12), .Q(\MEM[3] [30]), .QN());
   DFF_X1 \MEM_reg[3][29]  (.D(n_32_45), .CK(n_32_12), .Q(\MEM[3] [29]), .QN());
   DFF_X1 \MEM_reg[3][28]  (.D(n_32_44), .CK(n_32_12), .Q(\MEM[3] [28]), .QN());
   DFF_X1 \MEM_reg[3][27]  (.D(n_32_43), .CK(n_32_12), .Q(\MEM[3] [27]), .QN());
   DFF_X1 \MEM_reg[3][26]  (.D(n_32_42), .CK(n_32_12), .Q(\MEM[3] [26]), .QN());
   DFF_X1 \MEM_reg[3][25]  (.D(n_32_41), .CK(n_32_12), .Q(\MEM[3] [25]), .QN());
   DFF_X1 \MEM_reg[3][24]  (.D(n_32_40), .CK(n_32_12), .Q(\MEM[3] [24]), .QN());
   DFF_X1 \MEM_reg[3][23]  (.D(n_32_39), .CK(n_32_12), .Q(\MEM[3] [23]), .QN());
   DFF_X1 \MEM_reg[3][22]  (.D(n_32_38), .CK(n_32_12), .Q(\MEM[3] [22]), .QN());
   DFF_X1 \MEM_reg[3][21]  (.D(n_32_37), .CK(n_32_12), .Q(\MEM[3] [21]), .QN());
   DFF_X1 \MEM_reg[3][20]  (.D(n_32_36), .CK(n_32_12), .Q(\MEM[3] [20]), .QN());
   DFF_X1 \MEM_reg[3][19]  (.D(n_32_35), .CK(n_32_12), .Q(\MEM[3] [19]), .QN());
   DFF_X1 \MEM_reg[3][18]  (.D(n_32_34), .CK(n_32_12), .Q(\MEM[3] [18]), .QN());
   DFF_X1 \MEM_reg[3][17]  (.D(n_32_33), .CK(n_32_12), .Q(\MEM[3] [17]), .QN());
   DFF_X1 \MEM_reg[3][16]  (.D(n_32_32), .CK(n_32_12), .Q(\MEM[3] [16]), .QN());
   DFF_X1 \MEM_reg[3][15]  (.D(n_32_31), .CK(n_32_12), .Q(\MEM[3] [15]), .QN());
   DFF_X1 \MEM_reg[3][14]  (.D(n_32_30), .CK(n_32_12), .Q(\MEM[3] [14]), .QN());
   DFF_X1 \MEM_reg[3][13]  (.D(n_32_29), .CK(n_32_12), .Q(\MEM[3] [13]), .QN());
   DFF_X1 \MEM_reg[3][12]  (.D(n_32_28), .CK(n_32_12), .Q(\MEM[3] [12]), .QN());
   DFF_X1 \MEM_reg[3][11]  (.D(n_32_27), .CK(n_32_12), .Q(\MEM[3] [11]), .QN());
   DFF_X1 \MEM_reg[3][10]  (.D(n_32_26), .CK(n_32_12), .Q(\MEM[3] [10]), .QN());
   DFF_X1 \MEM_reg[3][9]  (.D(n_32_25), .CK(n_32_12), .Q(\MEM[3] [9]), .QN());
   DFF_X1 \MEM_reg[3][8]  (.D(n_32_24), .CK(n_32_12), .Q(\MEM[3] [8]), .QN());
   DFF_X1 \MEM_reg[3][7]  (.D(n_32_23), .CK(n_32_12), .Q(\MEM[3] [7]), .QN());
   DFF_X1 \MEM_reg[3][6]  (.D(n_32_22), .CK(n_32_12), .Q(\MEM[3] [6]), .QN());
   DFF_X1 \MEM_reg[3][5]  (.D(n_32_21), .CK(n_32_12), .Q(\MEM[3] [5]), .QN());
   DFF_X1 \MEM_reg[3][4]  (.D(n_32_20), .CK(n_32_12), .Q(\MEM[3] [4]), .QN());
   DFF_X1 \MEM_reg[3][3]  (.D(n_32_19), .CK(n_32_12), .Q(\MEM[3] [3]), .QN());
   DFF_X1 \MEM_reg[3][2]  (.D(n_32_18), .CK(n_32_12), .Q(\MEM[3] [2]), .QN());
   DFF_X1 \MEM_reg[3][1]  (.D(n_32_17), .CK(n_32_12), .Q(\MEM[3] [1]), .QN());
   DFF_X1 \MEM_reg[3][0]  (.D(n_32_16), .CK(n_32_12), .Q(\MEM[3] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[2]_reg  (.CK(clk), .E(n_32_50), .SE(1'b0), 
      .GCK(n_32_13));
   DFF_X1 \MEM_reg[2][31]  (.D(n_32_47), .CK(n_32_13), .Q(\MEM[2] [31]), .QN());
   DFF_X1 \MEM_reg[2][30]  (.D(n_32_46), .CK(n_32_13), .Q(\MEM[2] [30]), .QN());
   DFF_X1 \MEM_reg[2][29]  (.D(n_32_45), .CK(n_32_13), .Q(\MEM[2] [29]), .QN());
   DFF_X1 \MEM_reg[2][28]  (.D(n_32_44), .CK(n_32_13), .Q(\MEM[2] [28]), .QN());
   DFF_X1 \MEM_reg[2][27]  (.D(n_32_43), .CK(n_32_13), .Q(\MEM[2] [27]), .QN());
   DFF_X1 \MEM_reg[2][26]  (.D(n_32_42), .CK(n_32_13), .Q(\MEM[2] [26]), .QN());
   DFF_X1 \MEM_reg[2][25]  (.D(n_32_41), .CK(n_32_13), .Q(\MEM[2] [25]), .QN());
   DFF_X1 \MEM_reg[2][24]  (.D(n_32_40), .CK(n_32_13), .Q(\MEM[2] [24]), .QN());
   DFF_X1 \MEM_reg[2][23]  (.D(n_32_39), .CK(n_32_13), .Q(\MEM[2] [23]), .QN());
   DFF_X1 \MEM_reg[2][22]  (.D(n_32_38), .CK(n_32_13), .Q(\MEM[2] [22]), .QN());
   DFF_X1 \MEM_reg[2][21]  (.D(n_32_37), .CK(n_32_13), .Q(\MEM[2] [21]), .QN());
   DFF_X1 \MEM_reg[2][20]  (.D(n_32_36), .CK(n_32_13), .Q(\MEM[2] [20]), .QN());
   DFF_X1 \MEM_reg[2][19]  (.D(n_32_35), .CK(n_32_13), .Q(\MEM[2] [19]), .QN());
   DFF_X1 \MEM_reg[2][18]  (.D(n_32_34), .CK(n_32_13), .Q(\MEM[2] [18]), .QN());
   DFF_X1 \MEM_reg[2][17]  (.D(n_32_33), .CK(n_32_13), .Q(\MEM[2] [17]), .QN());
   DFF_X1 \MEM_reg[2][16]  (.D(n_32_32), .CK(n_32_13), .Q(\MEM[2] [16]), .QN());
   DFF_X1 \MEM_reg[2][15]  (.D(n_32_31), .CK(n_32_13), .Q(\MEM[2] [15]), .QN());
   DFF_X1 \MEM_reg[2][14]  (.D(n_32_30), .CK(n_32_13), .Q(\MEM[2] [14]), .QN());
   DFF_X1 \MEM_reg[2][13]  (.D(n_32_29), .CK(n_32_13), .Q(\MEM[2] [13]), .QN());
   DFF_X1 \MEM_reg[2][12]  (.D(n_32_28), .CK(n_32_13), .Q(\MEM[2] [12]), .QN());
   DFF_X1 \MEM_reg[2][11]  (.D(n_32_27), .CK(n_32_13), .Q(\MEM[2] [11]), .QN());
   DFF_X1 \MEM_reg[2][10]  (.D(n_32_26), .CK(n_32_13), .Q(\MEM[2] [10]), .QN());
   DFF_X1 \MEM_reg[2][9]  (.D(n_32_25), .CK(n_32_13), .Q(\MEM[2] [9]), .QN());
   DFF_X1 \MEM_reg[2][8]  (.D(n_32_24), .CK(n_32_13), .Q(\MEM[2] [8]), .QN());
   DFF_X1 \MEM_reg[2][7]  (.D(n_32_23), .CK(n_32_13), .Q(\MEM[2] [7]), .QN());
   DFF_X1 \MEM_reg[2][6]  (.D(n_32_22), .CK(n_32_13), .Q(\MEM[2] [6]), .QN());
   DFF_X1 \MEM_reg[2][5]  (.D(n_32_21), .CK(n_32_13), .Q(\MEM[2] [5]), .QN());
   DFF_X1 \MEM_reg[2][4]  (.D(n_32_20), .CK(n_32_13), .Q(\MEM[2] [4]), .QN());
   DFF_X1 \MEM_reg[2][3]  (.D(n_32_19), .CK(n_32_13), .Q(\MEM[2] [3]), .QN());
   DFF_X1 \MEM_reg[2][2]  (.D(n_32_18), .CK(n_32_13), .Q(\MEM[2] [2]), .QN());
   DFF_X1 \MEM_reg[2][1]  (.D(n_32_17), .CK(n_32_13), .Q(\MEM[2] [1]), .QN());
   DFF_X1 \MEM_reg[2][0]  (.D(n_32_16), .CK(n_32_13), .Q(\MEM[2] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[1]_reg  (.CK(clk), .E(n_32_49), .SE(1'b0), 
      .GCK(n_32_14));
   DFF_X1 \MEM_reg[1][31]  (.D(n_32_47), .CK(n_32_14), .Q(\MEM[1] [31]), .QN());
   DFF_X1 \MEM_reg[1][30]  (.D(n_32_46), .CK(n_32_14), .Q(\MEM[1] [30]), .QN());
   DFF_X1 \MEM_reg[1][29]  (.D(n_32_45), .CK(n_32_14), .Q(\MEM[1] [29]), .QN());
   DFF_X1 \MEM_reg[1][28]  (.D(n_32_44), .CK(n_32_14), .Q(\MEM[1] [28]), .QN());
   DFF_X1 \MEM_reg[1][27]  (.D(n_32_43), .CK(n_32_14), .Q(\MEM[1] [27]), .QN());
   DFF_X1 \MEM_reg[1][26]  (.D(n_32_42), .CK(n_32_14), .Q(\MEM[1] [26]), .QN());
   DFF_X1 \MEM_reg[1][25]  (.D(n_32_41), .CK(n_32_14), .Q(\MEM[1] [25]), .QN());
   DFF_X1 \MEM_reg[1][24]  (.D(n_32_40), .CK(n_32_14), .Q(\MEM[1] [24]), .QN());
   DFF_X1 \MEM_reg[1][23]  (.D(n_32_39), .CK(n_32_14), .Q(\MEM[1] [23]), .QN());
   DFF_X1 \MEM_reg[1][22]  (.D(n_32_38), .CK(n_32_14), .Q(\MEM[1] [22]), .QN());
   DFF_X1 \MEM_reg[1][21]  (.D(n_32_37), .CK(n_32_14), .Q(\MEM[1] [21]), .QN());
   DFF_X1 \MEM_reg[1][20]  (.D(n_32_36), .CK(n_32_14), .Q(\MEM[1] [20]), .QN());
   DFF_X1 \MEM_reg[1][19]  (.D(n_32_35), .CK(n_32_14), .Q(\MEM[1] [19]), .QN());
   DFF_X1 \MEM_reg[1][18]  (.D(n_32_34), .CK(n_32_14), .Q(\MEM[1] [18]), .QN());
   DFF_X1 \MEM_reg[1][17]  (.D(n_32_33), .CK(n_32_14), .Q(\MEM[1] [17]), .QN());
   DFF_X1 \MEM_reg[1][16]  (.D(n_32_32), .CK(n_32_14), .Q(\MEM[1] [16]), .QN());
   DFF_X1 \MEM_reg[1][15]  (.D(n_32_31), .CK(n_32_14), .Q(\MEM[1] [15]), .QN());
   DFF_X1 \MEM_reg[1][14]  (.D(n_32_30), .CK(n_32_14), .Q(\MEM[1] [14]), .QN());
   DFF_X1 \MEM_reg[1][13]  (.D(n_32_29), .CK(n_32_14), .Q(\MEM[1] [13]), .QN());
   DFF_X1 \MEM_reg[1][12]  (.D(n_32_28), .CK(n_32_14), .Q(\MEM[1] [12]), .QN());
   DFF_X1 \MEM_reg[1][11]  (.D(n_32_27), .CK(n_32_14), .Q(\MEM[1] [11]), .QN());
   DFF_X1 \MEM_reg[1][10]  (.D(n_32_26), .CK(n_32_14), .Q(\MEM[1] [10]), .QN());
   DFF_X1 \MEM_reg[1][9]  (.D(n_32_25), .CK(n_32_14), .Q(\MEM[1] [9]), .QN());
   DFF_X1 \MEM_reg[1][8]  (.D(n_32_24), .CK(n_32_14), .Q(\MEM[1] [8]), .QN());
   DFF_X1 \MEM_reg[1][7]  (.D(n_32_23), .CK(n_32_14), .Q(\MEM[1] [7]), .QN());
   DFF_X1 \MEM_reg[1][6]  (.D(n_32_22), .CK(n_32_14), .Q(\MEM[1] [6]), .QN());
   DFF_X1 \MEM_reg[1][5]  (.D(n_32_21), .CK(n_32_14), .Q(\MEM[1] [5]), .QN());
   DFF_X1 \MEM_reg[1][4]  (.D(n_32_20), .CK(n_32_14), .Q(\MEM[1] [4]), .QN());
   DFF_X1 \MEM_reg[1][3]  (.D(n_32_19), .CK(n_32_14), .Q(\MEM[1] [3]), .QN());
   DFF_X1 \MEM_reg[1][2]  (.D(n_32_18), .CK(n_32_14), .Q(\MEM[1] [2]), .QN());
   DFF_X1 \MEM_reg[1][1]  (.D(n_32_17), .CK(n_32_14), .Q(\MEM[1] [1]), .QN());
   DFF_X1 \MEM_reg[1][0]  (.D(n_32_16), .CK(n_32_14), .Q(\MEM[1] [0]), .QN());
   CLKGATETST_X1 \clk_gate_MEM_reg[0]_reg  (.CK(clk), .E(n_32_48), .SE(1'b0), 
      .GCK(n_32_15));
   DFF_X1 \MEM_reg[0][31]  (.D(n_32_47), .CK(n_32_15), .Q(\MEM[0] [31]), .QN());
   DFF_X1 \MEM_reg[0][30]  (.D(n_32_46), .CK(n_32_15), .Q(\MEM[0] [30]), .QN());
   DFF_X1 \MEM_reg[0][29]  (.D(n_32_45), .CK(n_32_15), .Q(\MEM[0] [29]), .QN());
   DFF_X1 \MEM_reg[0][28]  (.D(n_32_44), .CK(n_32_15), .Q(\MEM[0] [28]), .QN());
   DFF_X1 \MEM_reg[0][27]  (.D(n_32_43), .CK(n_32_15), .Q(\MEM[0] [27]), .QN());
   DFF_X1 \MEM_reg[0][26]  (.D(n_32_42), .CK(n_32_15), .Q(\MEM[0] [26]), .QN());
   DFF_X1 \MEM_reg[0][25]  (.D(n_32_41), .CK(n_32_15), .Q(\MEM[0] [25]), .QN());
   DFF_X1 \MEM_reg[0][24]  (.D(n_32_40), .CK(n_32_15), .Q(\MEM[0] [24]), .QN());
   DFF_X1 \MEM_reg[0][23]  (.D(n_32_39), .CK(n_32_15), .Q(\MEM[0] [23]), .QN());
   DFF_X1 \MEM_reg[0][22]  (.D(n_32_38), .CK(n_32_15), .Q(\MEM[0] [22]), .QN());
   DFF_X1 \MEM_reg[0][21]  (.D(n_32_37), .CK(n_32_15), .Q(\MEM[0] [21]), .QN());
   DFF_X1 \MEM_reg[0][20]  (.D(n_32_36), .CK(n_32_15), .Q(\MEM[0] [20]), .QN());
   DFF_X1 \MEM_reg[0][19]  (.D(n_32_35), .CK(n_32_15), .Q(\MEM[0] [19]), .QN());
   DFF_X1 \MEM_reg[0][18]  (.D(n_32_34), .CK(n_32_15), .Q(\MEM[0] [18]), .QN());
   DFF_X1 \MEM_reg[0][17]  (.D(n_32_33), .CK(n_32_15), .Q(\MEM[0] [17]), .QN());
   DFF_X1 \MEM_reg[0][16]  (.D(n_32_32), .CK(n_32_15), .Q(\MEM[0] [16]), .QN());
   DFF_X1 \MEM_reg[0][15]  (.D(n_32_31), .CK(n_32_15), .Q(\MEM[0] [15]), .QN());
   DFF_X1 \MEM_reg[0][14]  (.D(n_32_30), .CK(n_32_15), .Q(\MEM[0] [14]), .QN());
   DFF_X1 \MEM_reg[0][13]  (.D(n_32_29), .CK(n_32_15), .Q(\MEM[0] [13]), .QN());
   DFF_X1 \MEM_reg[0][12]  (.D(n_32_28), .CK(n_32_15), .Q(\MEM[0] [12]), .QN());
   DFF_X1 \MEM_reg[0][11]  (.D(n_32_27), .CK(n_32_15), .Q(\MEM[0] [11]), .QN());
   DFF_X1 \MEM_reg[0][10]  (.D(n_32_26), .CK(n_32_15), .Q(\MEM[0] [10]), .QN());
   DFF_X1 \MEM_reg[0][9]  (.D(n_32_25), .CK(n_32_15), .Q(\MEM[0] [9]), .QN());
   DFF_X1 \MEM_reg[0][8]  (.D(n_32_24), .CK(n_32_15), .Q(\MEM[0] [8]), .QN());
   DFF_X1 \MEM_reg[0][7]  (.D(n_32_23), .CK(n_32_15), .Q(\MEM[0] [7]), .QN());
   DFF_X1 \MEM_reg[0][6]  (.D(n_32_22), .CK(n_32_15), .Q(\MEM[0] [6]), .QN());
   DFF_X1 \MEM_reg[0][5]  (.D(n_32_21), .CK(n_32_15), .Q(\MEM[0] [5]), .QN());
   DFF_X1 \MEM_reg[0][4]  (.D(n_32_20), .CK(n_32_15), .Q(\MEM[0] [4]), .QN());
   DFF_X1 \MEM_reg[0][3]  (.D(n_32_19), .CK(n_32_15), .Q(\MEM[0] [3]), .QN());
   DFF_X1 \MEM_reg[0][2]  (.D(n_32_18), .CK(n_32_15), .Q(\MEM[0] [2]), .QN());
   DFF_X1 \MEM_reg[0][1]  (.D(n_32_17), .CK(n_32_15), .Q(\MEM[0] [1]), .QN());
   DFF_X1 \MEM_reg[0][0]  (.D(n_32_16), .CK(n_32_15), .Q(\MEM[0] [0]), .QN());
   INV_X1 i_32_0_0 (.A(addr1[0]), .ZN(n_32_0_0));
   OR2_X1 i_32_0_1 (.A1(n_32_0_0), .A2(addr1[1]), .ZN(n_32_0_1));
   INV_X1 i_32_0_2 (.A(addr1[2]), .ZN(n_32_0_2));
   NAND2_X1 i_32_0_3 (.A1(n_32_0_2), .A2(addr1[3]), .ZN(n_32_0_3));
   NOR2_X1 i_32_0_4 (.A1(n_32_0_1), .A2(n_32_0_3), .ZN(n_32_0_4));
   NAND2_X1 i_32_0_5 (.A1(n_32_0_0), .A2(addr1[1]), .ZN(n_32_0_5));
   NOR2_X1 i_32_0_6 (.A1(n_32_0_5), .A2(n_32_0_3), .ZN(n_32_0_6));
   AOI22_X1 i_32_0_7 (.A1(n_32_0_4), .A2(\MEM[9] [0]), .B1(n_32_0_6), .B2(
      \MEM[10] [0]), .ZN(n_32_0_7));
   OR2_X1 i_32_0_8 (.A1(n_32_0_2), .A2(addr1[3]), .ZN(n_32_0_8));
   NOR2_X1 i_32_0_9 (.A1(n_32_0_1), .A2(n_32_0_8), .ZN(n_32_0_9));
   OR2_X1 i_32_0_10 (.A1(addr1[3]), .A2(addr1[2]), .ZN(n_32_0_10));
   NAND2_X1 i_32_0_11 (.A1(addr1[0]), .A2(addr1[1]), .ZN(n_32_0_11));
   NOR2_X1 i_32_0_12 (.A1(n_32_0_10), .A2(n_32_0_11), .ZN(n_32_0_12));
   AOI22_X1 i_32_0_13 (.A1(n_32_0_9), .A2(\MEM[5] [0]), .B1(n_32_0_12), .B2(
      \MEM[3] [0]), .ZN(n_32_0_13));
   NOR2_X1 i_32_0_14 (.A1(n_32_0_8), .A2(n_32_0_5), .ZN(n_32_0_14));
   NOR2_X1 i_32_0_15 (.A1(n_32_0_8), .A2(n_32_0_11), .ZN(n_32_0_15));
   AOI22_X1 i_32_0_16 (.A1(\MEM[6] [0]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [0]), .ZN(n_32_0_16));
   OR2_X1 i_32_0_17 (.A1(addr1[0]), .A2(addr1[1]), .ZN(n_32_0_17));
   NOR2_X1 i_32_0_18 (.A1(n_32_0_17), .A2(n_32_0_3), .ZN(n_32_0_18));
   NOR2_X1 i_32_0_19 (.A1(n_32_0_3), .A2(n_32_0_11), .ZN(n_32_0_19));
   AOI22_X1 i_32_0_20 (.A1(\MEM[8] [0]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [0]), .ZN(n_32_0_20));
   NAND4_X1 i_32_0_21 (.A1(n_32_0_7), .A2(n_32_0_13), .A3(n_32_0_16), .A4(
      n_32_0_20), .ZN(n_32_0_21));
   NOR2_X1 i_32_0_22 (.A1(n_32_0_10), .A2(n_32_0_5), .ZN(n_32_0_22));
   NOR2_X1 i_32_0_23 (.A1(n_32_0_17), .A2(n_32_0_10), .ZN(n_32_0_23));
   AOI221_X1 i_32_0_24 (.A(n_32_0_21), .B1(\MEM[2] [0]), .B2(n_32_0_22), 
      .C1(\MEM[0] [0]), .C2(n_32_0_23), .ZN(n_32_0_24));
   NOR2_X1 i_32_0_25 (.A1(n_32_0_8), .A2(n_32_0_17), .ZN(n_32_0_25));
   NAND2_X1 i_32_0_26 (.A1(addr1[3]), .A2(addr1[2]), .ZN(n_32_0_26));
   NOR2_X1 i_32_0_27 (.A1(n_32_0_1), .A2(n_32_0_26), .ZN(n_32_0_27));
   AOI22_X1 i_32_0_28 (.A1(\MEM[4] [0]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [0]), .ZN(n_32_0_28));
   NOR2_X1 i_32_0_29 (.A1(n_32_0_1), .A2(n_32_0_10), .ZN(n_32_0_29));
   NOR2_X1 i_32_0_30 (.A1(n_32_0_26), .A2(n_32_0_11), .ZN(n_32_0_30));
   AOI22_X1 i_32_0_31 (.A1(\MEM[1] [0]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [0]), .ZN(n_32_0_31));
   NOR2_X1 i_32_0_32 (.A1(n_32_0_17), .A2(n_32_0_26), .ZN(n_32_0_32));
   NOR2_X1 i_32_0_33 (.A1(n_32_0_5), .A2(n_32_0_26), .ZN(n_32_0_33));
   AOI22_X1 i_32_0_34 (.A1(\MEM[12] [0]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [0]), .ZN(n_32_0_34));
   NAND4_X1 i_32_0_35 (.A1(n_32_0_24), .A2(n_32_0_28), .A3(n_32_0_31), .A4(
      n_32_0_34), .ZN(MEM[0]));
   INV_X1 i_32_0_36 (.A(we1), .ZN(n_32_0_35));
   OAI22_X1 i_32_0_37 (.A1(MEM[0]), .A2(we1), .B1(data1[0]), .B2(n_32_0_35), 
      .ZN(n_32_0_36));
   NOR2_X1 i_32_0_38 (.A1(n_32_0_36), .A2(rst), .ZN(n_32_16));
   AOI22_X1 i_32_0_39 (.A1(n_32_0_4), .A2(\MEM[9] [1]), .B1(n_32_0_6), .B2(
      \MEM[10] [1]), .ZN(n_32_0_37));
   AOI22_X1 i_32_0_40 (.A1(n_32_0_9), .A2(\MEM[5] [1]), .B1(n_32_0_12), .B2(
      \MEM[3] [1]), .ZN(n_32_0_38));
   AOI22_X1 i_32_0_41 (.A1(\MEM[6] [1]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [1]), .ZN(n_32_0_39));
   AOI22_X1 i_32_0_42 (.A1(\MEM[8] [1]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [1]), .ZN(n_32_0_40));
   NAND4_X1 i_32_0_43 (.A1(n_32_0_37), .A2(n_32_0_38), .A3(n_32_0_39), .A4(
      n_32_0_40), .ZN(n_32_0_41));
   AOI221_X1 i_32_0_44 (.A(n_32_0_41), .B1(\MEM[2] [1]), .B2(n_32_0_22), 
      .C1(\MEM[0] [1]), .C2(n_32_0_23), .ZN(n_32_0_42));
   AOI22_X1 i_32_0_45 (.A1(\MEM[4] [1]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [1]), .ZN(n_32_0_43));
   AOI22_X1 i_32_0_46 (.A1(\MEM[1] [1]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [1]), .ZN(n_32_0_44));
   AOI22_X1 i_32_0_47 (.A1(\MEM[12] [1]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [1]), .ZN(n_32_0_45));
   NAND4_X1 i_32_0_48 (.A1(n_32_0_42), .A2(n_32_0_43), .A3(n_32_0_44), .A4(
      n_32_0_45), .ZN(MEM[1]));
   OAI22_X1 i_32_0_49 (.A1(MEM[1]), .A2(we1), .B1(data1[1]), .B2(n_32_0_35), 
      .ZN(n_32_0_46));
   NOR2_X1 i_32_0_50 (.A1(n_32_0_46), .A2(rst), .ZN(n_32_17));
   AOI22_X1 i_32_0_51 (.A1(n_32_0_4), .A2(\MEM[9] [2]), .B1(n_32_0_6), .B2(
      \MEM[10] [2]), .ZN(n_32_0_47));
   AOI22_X1 i_32_0_52 (.A1(n_32_0_9), .A2(\MEM[5] [2]), .B1(n_32_0_12), .B2(
      \MEM[3] [2]), .ZN(n_32_0_48));
   AOI22_X1 i_32_0_53 (.A1(\MEM[6] [2]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [2]), .ZN(n_32_0_49));
   AOI22_X1 i_32_0_54 (.A1(\MEM[8] [2]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [2]), .ZN(n_32_0_50));
   NAND4_X1 i_32_0_55 (.A1(n_32_0_47), .A2(n_32_0_48), .A3(n_32_0_49), .A4(
      n_32_0_50), .ZN(n_32_0_51));
   AOI221_X1 i_32_0_56 (.A(n_32_0_51), .B1(\MEM[2] [2]), .B2(n_32_0_22), 
      .C1(\MEM[0] [2]), .C2(n_32_0_23), .ZN(n_32_0_52));
   AOI22_X1 i_32_0_57 (.A1(\MEM[4] [2]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [2]), .ZN(n_32_0_53));
   AOI22_X1 i_32_0_58 (.A1(\MEM[1] [2]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [2]), .ZN(n_32_0_54));
   AOI22_X1 i_32_0_59 (.A1(\MEM[12] [2]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [2]), .ZN(n_32_0_55));
   NAND4_X1 i_32_0_60 (.A1(n_32_0_52), .A2(n_32_0_53), .A3(n_32_0_54), .A4(
      n_32_0_55), .ZN(MEM[2]));
   OAI22_X1 i_32_0_61 (.A1(MEM[2]), .A2(we1), .B1(data1[2]), .B2(n_32_0_35), 
      .ZN(n_32_0_56));
   NOR2_X1 i_32_0_62 (.A1(n_32_0_56), .A2(rst), .ZN(n_32_18));
   AOI22_X1 i_32_0_63 (.A1(n_32_0_4), .A2(\MEM[9] [3]), .B1(n_32_0_6), .B2(
      \MEM[10] [3]), .ZN(n_32_0_57));
   AOI22_X1 i_32_0_64 (.A1(n_32_0_9), .A2(\MEM[5] [3]), .B1(n_32_0_12), .B2(
      \MEM[3] [3]), .ZN(n_32_0_58));
   AOI22_X1 i_32_0_65 (.A1(\MEM[6] [3]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [3]), .ZN(n_32_0_59));
   AOI22_X1 i_32_0_66 (.A1(\MEM[8] [3]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [3]), .ZN(n_32_0_60));
   NAND4_X1 i_32_0_67 (.A1(n_32_0_57), .A2(n_32_0_58), .A3(n_32_0_59), .A4(
      n_32_0_60), .ZN(n_32_0_61));
   AOI221_X1 i_32_0_68 (.A(n_32_0_61), .B1(\MEM[2] [3]), .B2(n_32_0_22), 
      .C1(\MEM[0] [3]), .C2(n_32_0_23), .ZN(n_32_0_62));
   AOI22_X1 i_32_0_69 (.A1(\MEM[4] [3]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [3]), .ZN(n_32_0_63));
   AOI22_X1 i_32_0_70 (.A1(\MEM[1] [3]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [3]), .ZN(n_32_0_64));
   AOI22_X1 i_32_0_71 (.A1(\MEM[12] [3]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [3]), .ZN(n_32_0_65));
   NAND4_X1 i_32_0_72 (.A1(n_32_0_62), .A2(n_32_0_63), .A3(n_32_0_64), .A4(
      n_32_0_65), .ZN(MEM[3]));
   OAI22_X1 i_32_0_73 (.A1(MEM[3]), .A2(we1), .B1(data1[3]), .B2(n_32_0_35), 
      .ZN(n_32_0_66));
   NOR2_X1 i_32_0_74 (.A1(n_32_0_66), .A2(rst), .ZN(n_32_19));
   AOI22_X1 i_32_0_75 (.A1(n_32_0_4), .A2(\MEM[9] [4]), .B1(n_32_0_6), .B2(
      \MEM[10] [4]), .ZN(n_32_0_67));
   AOI22_X1 i_32_0_76 (.A1(n_32_0_9), .A2(\MEM[5] [4]), .B1(n_32_0_12), .B2(
      \MEM[3] [4]), .ZN(n_32_0_68));
   AOI22_X1 i_32_0_77 (.A1(\MEM[6] [4]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [4]), .ZN(n_32_0_69));
   AOI22_X1 i_32_0_78 (.A1(\MEM[8] [4]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [4]), .ZN(n_32_0_70));
   NAND4_X1 i_32_0_79 (.A1(n_32_0_67), .A2(n_32_0_68), .A3(n_32_0_69), .A4(
      n_32_0_70), .ZN(n_32_0_71));
   AOI221_X1 i_32_0_80 (.A(n_32_0_71), .B1(\MEM[2] [4]), .B2(n_32_0_22), 
      .C1(\MEM[0] [4]), .C2(n_32_0_23), .ZN(n_32_0_72));
   AOI22_X1 i_32_0_81 (.A1(\MEM[4] [4]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [4]), .ZN(n_32_0_73));
   AOI22_X1 i_32_0_82 (.A1(\MEM[1] [4]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [4]), .ZN(n_32_0_74));
   AOI22_X1 i_32_0_83 (.A1(\MEM[12] [4]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [4]), .ZN(n_32_0_75));
   NAND4_X1 i_32_0_84 (.A1(n_32_0_72), .A2(n_32_0_73), .A3(n_32_0_74), .A4(
      n_32_0_75), .ZN(MEM[4]));
   OAI22_X1 i_32_0_85 (.A1(MEM[4]), .A2(we1), .B1(data1[4]), .B2(n_32_0_35), 
      .ZN(n_32_0_76));
   NOR2_X1 i_32_0_86 (.A1(n_32_0_76), .A2(rst), .ZN(n_32_20));
   AOI22_X1 i_32_0_87 (.A1(n_32_0_4), .A2(\MEM[9] [5]), .B1(n_32_0_6), .B2(
      \MEM[10] [5]), .ZN(n_32_0_77));
   AOI22_X1 i_32_0_88 (.A1(n_32_0_9), .A2(\MEM[5] [5]), .B1(n_32_0_12), .B2(
      \MEM[3] [5]), .ZN(n_32_0_78));
   AOI22_X1 i_32_0_89 (.A1(\MEM[6] [5]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [5]), .ZN(n_32_0_79));
   AOI22_X1 i_32_0_90 (.A1(\MEM[8] [5]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [5]), .ZN(n_32_0_80));
   NAND4_X1 i_32_0_91 (.A1(n_32_0_77), .A2(n_32_0_78), .A3(n_32_0_79), .A4(
      n_32_0_80), .ZN(n_32_0_81));
   AOI221_X1 i_32_0_92 (.A(n_32_0_81), .B1(\MEM[2] [5]), .B2(n_32_0_22), 
      .C1(\MEM[0] [5]), .C2(n_32_0_23), .ZN(n_32_0_82));
   AOI22_X1 i_32_0_93 (.A1(\MEM[4] [5]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [5]), .ZN(n_32_0_83));
   AOI22_X1 i_32_0_94 (.A1(\MEM[1] [5]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [5]), .ZN(n_32_0_84));
   AOI22_X1 i_32_0_95 (.A1(\MEM[12] [5]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [5]), .ZN(n_32_0_85));
   NAND4_X1 i_32_0_96 (.A1(n_32_0_82), .A2(n_32_0_83), .A3(n_32_0_84), .A4(
      n_32_0_85), .ZN(MEM[5]));
   OAI22_X1 i_32_0_97 (.A1(MEM[5]), .A2(we1), .B1(data1[5]), .B2(n_32_0_35), 
      .ZN(n_32_0_86));
   NOR2_X1 i_32_0_98 (.A1(n_32_0_86), .A2(rst), .ZN(n_32_21));
   AOI22_X1 i_32_0_99 (.A1(n_32_0_4), .A2(\MEM[9] [6]), .B1(n_32_0_6), .B2(
      \MEM[10] [6]), .ZN(n_32_0_87));
   AOI22_X1 i_32_0_100 (.A1(n_32_0_9), .A2(\MEM[5] [6]), .B1(n_32_0_12), 
      .B2(\MEM[3] [6]), .ZN(n_32_0_88));
   AOI22_X1 i_32_0_101 (.A1(\MEM[6] [6]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [6]), .ZN(n_32_0_89));
   AOI22_X1 i_32_0_102 (.A1(\MEM[8] [6]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [6]), .ZN(n_32_0_90));
   NAND4_X1 i_32_0_103 (.A1(n_32_0_87), .A2(n_32_0_88), .A3(n_32_0_89), .A4(
      n_32_0_90), .ZN(n_32_0_91));
   AOI221_X1 i_32_0_104 (.A(n_32_0_91), .B1(\MEM[2] [6]), .B2(n_32_0_22), 
      .C1(\MEM[0] [6]), .C2(n_32_0_23), .ZN(n_32_0_92));
   AOI22_X1 i_32_0_105 (.A1(\MEM[4] [6]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [6]), .ZN(n_32_0_93));
   AOI22_X1 i_32_0_106 (.A1(\MEM[1] [6]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [6]), .ZN(n_32_0_94));
   AOI22_X1 i_32_0_107 (.A1(\MEM[12] [6]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [6]), .ZN(n_32_0_95));
   NAND4_X1 i_32_0_108 (.A1(n_32_0_92), .A2(n_32_0_93), .A3(n_32_0_94), .A4(
      n_32_0_95), .ZN(MEM[6]));
   OAI22_X1 i_32_0_109 (.A1(MEM[6]), .A2(we1), .B1(data1[6]), .B2(n_32_0_35), 
      .ZN(n_32_0_96));
   NOR2_X1 i_32_0_110 (.A1(n_32_0_96), .A2(rst), .ZN(n_32_22));
   AOI22_X1 i_32_0_111 (.A1(n_32_0_4), .A2(\MEM[9] [7]), .B1(n_32_0_6), .B2(
      \MEM[10] [7]), .ZN(n_32_0_97));
   AOI22_X1 i_32_0_112 (.A1(n_32_0_9), .A2(\MEM[5] [7]), .B1(n_32_0_12), 
      .B2(\MEM[3] [7]), .ZN(n_32_0_98));
   AOI22_X1 i_32_0_113 (.A1(\MEM[6] [7]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [7]), .ZN(n_32_0_99));
   AOI22_X1 i_32_0_114 (.A1(\MEM[8] [7]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [7]), .ZN(n_32_0_100));
   NAND4_X1 i_32_0_115 (.A1(n_32_0_97), .A2(n_32_0_98), .A3(n_32_0_99), .A4(
      n_32_0_100), .ZN(n_32_0_101));
   AOI221_X1 i_32_0_116 (.A(n_32_0_101), .B1(\MEM[2] [7]), .B2(n_32_0_22), 
      .C1(\MEM[0] [7]), .C2(n_32_0_23), .ZN(n_32_0_102));
   AOI22_X1 i_32_0_117 (.A1(\MEM[4] [7]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [7]), .ZN(n_32_0_103));
   AOI22_X1 i_32_0_118 (.A1(\MEM[1] [7]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [7]), .ZN(n_32_0_104));
   AOI22_X1 i_32_0_119 (.A1(\MEM[12] [7]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [7]), .ZN(n_32_0_105));
   NAND4_X1 i_32_0_120 (.A1(n_32_0_102), .A2(n_32_0_103), .A3(n_32_0_104), 
      .A4(n_32_0_105), .ZN(MEM[7]));
   OAI22_X1 i_32_0_121 (.A1(MEM[7]), .A2(we1), .B1(data1[7]), .B2(n_32_0_35), 
      .ZN(n_32_0_106));
   NOR2_X1 i_32_0_122 (.A1(n_32_0_106), .A2(rst), .ZN(n_32_23));
   AOI22_X1 i_32_0_123 (.A1(n_32_0_4), .A2(\MEM[9] [8]), .B1(n_32_0_6), .B2(
      \MEM[10] [8]), .ZN(n_32_0_107));
   AOI22_X1 i_32_0_124 (.A1(n_32_0_9), .A2(\MEM[5] [8]), .B1(n_32_0_12), 
      .B2(\MEM[3] [8]), .ZN(n_32_0_108));
   AOI22_X1 i_32_0_125 (.A1(\MEM[6] [8]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [8]), .ZN(n_32_0_109));
   AOI22_X1 i_32_0_126 (.A1(\MEM[8] [8]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [8]), .ZN(n_32_0_110));
   NAND4_X1 i_32_0_127 (.A1(n_32_0_107), .A2(n_32_0_108), .A3(n_32_0_109), 
      .A4(n_32_0_110), .ZN(n_32_0_111));
   AOI221_X1 i_32_0_128 (.A(n_32_0_111), .B1(\MEM[2] [8]), .B2(n_32_0_22), 
      .C1(\MEM[0] [8]), .C2(n_32_0_23), .ZN(n_32_0_112));
   AOI22_X1 i_32_0_129 (.A1(\MEM[4] [8]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [8]), .ZN(n_32_0_113));
   AOI22_X1 i_32_0_130 (.A1(\MEM[1] [8]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [8]), .ZN(n_32_0_114));
   AOI22_X1 i_32_0_131 (.A1(\MEM[12] [8]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [8]), .ZN(n_32_0_115));
   NAND4_X1 i_32_0_132 (.A1(n_32_0_112), .A2(n_32_0_113), .A3(n_32_0_114), 
      .A4(n_32_0_115), .ZN(MEM[8]));
   OAI22_X1 i_32_0_133 (.A1(MEM[8]), .A2(we1), .B1(data1[8]), .B2(n_32_0_35), 
      .ZN(n_32_0_116));
   NOR2_X1 i_32_0_134 (.A1(n_32_0_116), .A2(rst), .ZN(n_32_24));
   AOI22_X1 i_32_0_135 (.A1(n_32_0_4), .A2(\MEM[9] [9]), .B1(n_32_0_6), .B2(
      \MEM[10] [9]), .ZN(n_32_0_117));
   AOI22_X1 i_32_0_136 (.A1(n_32_0_9), .A2(\MEM[5] [9]), .B1(n_32_0_12), 
      .B2(\MEM[3] [9]), .ZN(n_32_0_118));
   AOI22_X1 i_32_0_137 (.A1(\MEM[6] [9]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [9]), .ZN(n_32_0_119));
   AOI22_X1 i_32_0_138 (.A1(\MEM[8] [9]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [9]), .ZN(n_32_0_120));
   NAND4_X1 i_32_0_139 (.A1(n_32_0_117), .A2(n_32_0_118), .A3(n_32_0_119), 
      .A4(n_32_0_120), .ZN(n_32_0_121));
   AOI221_X1 i_32_0_140 (.A(n_32_0_121), .B1(\MEM[2] [9]), .B2(n_32_0_22), 
      .C1(\MEM[0] [9]), .C2(n_32_0_23), .ZN(n_32_0_122));
   AOI22_X1 i_32_0_141 (.A1(\MEM[4] [9]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [9]), .ZN(n_32_0_123));
   AOI22_X1 i_32_0_142 (.A1(\MEM[1] [9]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [9]), .ZN(n_32_0_124));
   AOI22_X1 i_32_0_143 (.A1(\MEM[12] [9]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [9]), .ZN(n_32_0_125));
   NAND4_X1 i_32_0_144 (.A1(n_32_0_122), .A2(n_32_0_123), .A3(n_32_0_124), 
      .A4(n_32_0_125), .ZN(MEM[9]));
   OAI22_X1 i_32_0_145 (.A1(MEM[9]), .A2(we1), .B1(data1[9]), .B2(n_32_0_35), 
      .ZN(n_32_0_126));
   NOR2_X1 i_32_0_146 (.A1(n_32_0_126), .A2(rst), .ZN(n_32_25));
   AOI22_X1 i_32_0_147 (.A1(n_32_0_4), .A2(\MEM[9] [10]), .B1(n_32_0_6), 
      .B2(\MEM[10] [10]), .ZN(n_32_0_127));
   AOI22_X1 i_32_0_148 (.A1(n_32_0_9), .A2(\MEM[5] [10]), .B1(n_32_0_12), 
      .B2(\MEM[3] [10]), .ZN(n_32_0_128));
   AOI22_X1 i_32_0_149 (.A1(\MEM[6] [10]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [10]), .ZN(n_32_0_129));
   AOI22_X1 i_32_0_150 (.A1(\MEM[8] [10]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [10]), .ZN(n_32_0_130));
   NAND4_X1 i_32_0_151 (.A1(n_32_0_127), .A2(n_32_0_128), .A3(n_32_0_129), 
      .A4(n_32_0_130), .ZN(n_32_0_131));
   AOI221_X1 i_32_0_152 (.A(n_32_0_131), .B1(\MEM[2] [10]), .B2(n_32_0_22), 
      .C1(\MEM[0] [10]), .C2(n_32_0_23), .ZN(n_32_0_132));
   AOI22_X1 i_32_0_153 (.A1(\MEM[4] [10]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [10]), .ZN(n_32_0_133));
   AOI22_X1 i_32_0_154 (.A1(\MEM[1] [10]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [10]), .ZN(n_32_0_134));
   AOI22_X1 i_32_0_155 (.A1(\MEM[12] [10]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [10]), .ZN(n_32_0_135));
   NAND4_X1 i_32_0_156 (.A1(n_32_0_132), .A2(n_32_0_133), .A3(n_32_0_134), 
      .A4(n_32_0_135), .ZN(MEM[10]));
   OAI22_X1 i_32_0_157 (.A1(MEM[10]), .A2(we1), .B1(data1[10]), .B2(n_32_0_35), 
      .ZN(n_32_0_136));
   NOR2_X1 i_32_0_158 (.A1(n_32_0_136), .A2(rst), .ZN(n_32_26));
   AOI22_X1 i_32_0_159 (.A1(n_32_0_4), .A2(\MEM[9] [11]), .B1(n_32_0_6), 
      .B2(\MEM[10] [11]), .ZN(n_32_0_137));
   AOI22_X1 i_32_0_160 (.A1(n_32_0_9), .A2(\MEM[5] [11]), .B1(n_32_0_12), 
      .B2(\MEM[3] [11]), .ZN(n_32_0_138));
   AOI22_X1 i_32_0_161 (.A1(\MEM[6] [11]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [11]), .ZN(n_32_0_139));
   AOI22_X1 i_32_0_162 (.A1(\MEM[8] [11]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [11]), .ZN(n_32_0_140));
   NAND4_X1 i_32_0_163 (.A1(n_32_0_137), .A2(n_32_0_138), .A3(n_32_0_139), 
      .A4(n_32_0_140), .ZN(n_32_0_141));
   AOI221_X1 i_32_0_164 (.A(n_32_0_141), .B1(\MEM[2] [11]), .B2(n_32_0_22), 
      .C1(\MEM[0] [11]), .C2(n_32_0_23), .ZN(n_32_0_142));
   AOI22_X1 i_32_0_165 (.A1(\MEM[4] [11]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [11]), .ZN(n_32_0_143));
   AOI22_X1 i_32_0_166 (.A1(\MEM[1] [11]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [11]), .ZN(n_32_0_144));
   AOI22_X1 i_32_0_167 (.A1(\MEM[12] [11]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [11]), .ZN(n_32_0_145));
   NAND4_X1 i_32_0_168 (.A1(n_32_0_142), .A2(n_32_0_143), .A3(n_32_0_144), 
      .A4(n_32_0_145), .ZN(MEM[11]));
   OAI22_X1 i_32_0_169 (.A1(MEM[11]), .A2(we1), .B1(data1[11]), .B2(n_32_0_35), 
      .ZN(n_32_0_146));
   NOR2_X1 i_32_0_170 (.A1(n_32_0_146), .A2(rst), .ZN(n_32_27));
   AOI22_X1 i_32_0_171 (.A1(n_32_0_4), .A2(\MEM[9] [12]), .B1(n_32_0_6), 
      .B2(\MEM[10] [12]), .ZN(n_32_0_147));
   AOI22_X1 i_32_0_172 (.A1(n_32_0_9), .A2(\MEM[5] [12]), .B1(n_32_0_12), 
      .B2(\MEM[3] [12]), .ZN(n_32_0_148));
   AOI22_X1 i_32_0_173 (.A1(\MEM[6] [12]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [12]), .ZN(n_32_0_149));
   AOI22_X1 i_32_0_174 (.A1(\MEM[8] [12]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [12]), .ZN(n_32_0_150));
   NAND4_X1 i_32_0_175 (.A1(n_32_0_147), .A2(n_32_0_148), .A3(n_32_0_149), 
      .A4(n_32_0_150), .ZN(n_32_0_151));
   AOI221_X1 i_32_0_176 (.A(n_32_0_151), .B1(\MEM[2] [12]), .B2(n_32_0_22), 
      .C1(\MEM[0] [12]), .C2(n_32_0_23), .ZN(n_32_0_152));
   AOI22_X1 i_32_0_177 (.A1(\MEM[4] [12]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [12]), .ZN(n_32_0_153));
   AOI22_X1 i_32_0_178 (.A1(\MEM[1] [12]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [12]), .ZN(n_32_0_154));
   AOI22_X1 i_32_0_179 (.A1(\MEM[12] [12]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [12]), .ZN(n_32_0_155));
   NAND4_X1 i_32_0_180 (.A1(n_32_0_152), .A2(n_32_0_153), .A3(n_32_0_154), 
      .A4(n_32_0_155), .ZN(MEM[12]));
   OAI22_X1 i_32_0_181 (.A1(MEM[12]), .A2(we1), .B1(data1[12]), .B2(n_32_0_35), 
      .ZN(n_32_0_156));
   NOR2_X1 i_32_0_182 (.A1(n_32_0_156), .A2(rst), .ZN(n_32_28));
   AOI22_X1 i_32_0_183 (.A1(n_32_0_4), .A2(\MEM[9] [13]), .B1(n_32_0_6), 
      .B2(\MEM[10] [13]), .ZN(n_32_0_157));
   AOI22_X1 i_32_0_184 (.A1(n_32_0_9), .A2(\MEM[5] [13]), .B1(n_32_0_12), 
      .B2(\MEM[3] [13]), .ZN(n_32_0_158));
   AOI22_X1 i_32_0_185 (.A1(\MEM[6] [13]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [13]), .ZN(n_32_0_159));
   AOI22_X1 i_32_0_186 (.A1(\MEM[8] [13]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [13]), .ZN(n_32_0_160));
   NAND4_X1 i_32_0_187 (.A1(n_32_0_157), .A2(n_32_0_158), .A3(n_32_0_159), 
      .A4(n_32_0_160), .ZN(n_32_0_161));
   AOI221_X1 i_32_0_188 (.A(n_32_0_161), .B1(\MEM[2] [13]), .B2(n_32_0_22), 
      .C1(\MEM[0] [13]), .C2(n_32_0_23), .ZN(n_32_0_162));
   AOI22_X1 i_32_0_189 (.A1(\MEM[4] [13]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [13]), .ZN(n_32_0_163));
   AOI22_X1 i_32_0_190 (.A1(\MEM[1] [13]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [13]), .ZN(n_32_0_164));
   AOI22_X1 i_32_0_191 (.A1(\MEM[12] [13]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [13]), .ZN(n_32_0_165));
   NAND4_X1 i_32_0_192 (.A1(n_32_0_162), .A2(n_32_0_163), .A3(n_32_0_164), 
      .A4(n_32_0_165), .ZN(MEM[13]));
   OAI22_X1 i_32_0_193 (.A1(MEM[13]), .A2(we1), .B1(data1[13]), .B2(n_32_0_35), 
      .ZN(n_32_0_166));
   NOR2_X1 i_32_0_194 (.A1(n_32_0_166), .A2(rst), .ZN(n_32_29));
   AOI22_X1 i_32_0_195 (.A1(n_32_0_4), .A2(\MEM[9] [14]), .B1(n_32_0_6), 
      .B2(\MEM[10] [14]), .ZN(n_32_0_167));
   AOI22_X1 i_32_0_196 (.A1(n_32_0_9), .A2(\MEM[5] [14]), .B1(n_32_0_12), 
      .B2(\MEM[3] [14]), .ZN(n_32_0_168));
   AOI22_X1 i_32_0_197 (.A1(\MEM[6] [14]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [14]), .ZN(n_32_0_169));
   AOI22_X1 i_32_0_198 (.A1(\MEM[8] [14]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [14]), .ZN(n_32_0_170));
   NAND4_X1 i_32_0_199 (.A1(n_32_0_167), .A2(n_32_0_168), .A3(n_32_0_169), 
      .A4(n_32_0_170), .ZN(n_32_0_171));
   AOI221_X1 i_32_0_200 (.A(n_32_0_171), .B1(\MEM[2] [14]), .B2(n_32_0_22), 
      .C1(\MEM[0] [14]), .C2(n_32_0_23), .ZN(n_32_0_172));
   AOI22_X1 i_32_0_201 (.A1(\MEM[4] [14]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [14]), .ZN(n_32_0_173));
   AOI22_X1 i_32_0_202 (.A1(\MEM[1] [14]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [14]), .ZN(n_32_0_174));
   AOI22_X1 i_32_0_203 (.A1(\MEM[12] [14]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [14]), .ZN(n_32_0_175));
   NAND4_X1 i_32_0_204 (.A1(n_32_0_172), .A2(n_32_0_173), .A3(n_32_0_174), 
      .A4(n_32_0_175), .ZN(MEM[14]));
   OAI22_X1 i_32_0_205 (.A1(MEM[14]), .A2(we1), .B1(data1[14]), .B2(n_32_0_35), 
      .ZN(n_32_0_176));
   NOR2_X1 i_32_0_206 (.A1(n_32_0_176), .A2(rst), .ZN(n_32_30));
   AOI22_X1 i_32_0_207 (.A1(n_32_0_4), .A2(\MEM[9] [15]), .B1(n_32_0_6), 
      .B2(\MEM[10] [15]), .ZN(n_32_0_177));
   AOI22_X1 i_32_0_208 (.A1(n_32_0_9), .A2(\MEM[5] [15]), .B1(n_32_0_12), 
      .B2(\MEM[3] [15]), .ZN(n_32_0_178));
   AOI22_X1 i_32_0_209 (.A1(\MEM[6] [15]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [15]), .ZN(n_32_0_179));
   AOI22_X1 i_32_0_210 (.A1(\MEM[8] [15]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [15]), .ZN(n_32_0_180));
   NAND4_X1 i_32_0_211 (.A1(n_32_0_177), .A2(n_32_0_178), .A3(n_32_0_179), 
      .A4(n_32_0_180), .ZN(n_32_0_181));
   AOI221_X1 i_32_0_212 (.A(n_32_0_181), .B1(\MEM[2] [15]), .B2(n_32_0_22), 
      .C1(\MEM[0] [15]), .C2(n_32_0_23), .ZN(n_32_0_182));
   AOI22_X1 i_32_0_213 (.A1(\MEM[4] [15]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [15]), .ZN(n_32_0_183));
   AOI22_X1 i_32_0_214 (.A1(\MEM[1] [15]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [15]), .ZN(n_32_0_184));
   AOI22_X1 i_32_0_215 (.A1(\MEM[12] [15]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [15]), .ZN(n_32_0_185));
   NAND4_X1 i_32_0_216 (.A1(n_32_0_182), .A2(n_32_0_183), .A3(n_32_0_184), 
      .A4(n_32_0_185), .ZN(MEM[15]));
   OAI22_X1 i_32_0_217 (.A1(MEM[15]), .A2(we1), .B1(data1[15]), .B2(n_32_0_35), 
      .ZN(n_32_0_186));
   NOR2_X1 i_32_0_218 (.A1(n_32_0_186), .A2(rst), .ZN(n_32_31));
   AOI22_X1 i_32_0_219 (.A1(n_32_0_4), .A2(\MEM[9] [16]), .B1(n_32_0_6), 
      .B2(\MEM[10] [16]), .ZN(n_32_0_187));
   AOI22_X1 i_32_0_220 (.A1(n_32_0_9), .A2(\MEM[5] [16]), .B1(n_32_0_12), 
      .B2(\MEM[3] [16]), .ZN(n_32_0_188));
   AOI22_X1 i_32_0_221 (.A1(\MEM[6] [16]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [16]), .ZN(n_32_0_189));
   AOI22_X1 i_32_0_222 (.A1(\MEM[8] [16]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [16]), .ZN(n_32_0_190));
   NAND4_X1 i_32_0_223 (.A1(n_32_0_187), .A2(n_32_0_188), .A3(n_32_0_189), 
      .A4(n_32_0_190), .ZN(n_32_0_191));
   AOI221_X1 i_32_0_224 (.A(n_32_0_191), .B1(\MEM[2] [16]), .B2(n_32_0_22), 
      .C1(\MEM[0] [16]), .C2(n_32_0_23), .ZN(n_32_0_192));
   AOI22_X1 i_32_0_225 (.A1(\MEM[4] [16]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [16]), .ZN(n_32_0_193));
   AOI22_X1 i_32_0_226 (.A1(\MEM[1] [16]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [16]), .ZN(n_32_0_194));
   AOI22_X1 i_32_0_227 (.A1(\MEM[12] [16]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [16]), .ZN(n_32_0_195));
   NAND4_X1 i_32_0_228 (.A1(n_32_0_192), .A2(n_32_0_193), .A3(n_32_0_194), 
      .A4(n_32_0_195), .ZN(MEM[16]));
   OAI22_X1 i_32_0_229 (.A1(MEM[16]), .A2(we1), .B1(data1[16]), .B2(n_32_0_35), 
      .ZN(n_32_0_196));
   NOR2_X1 i_32_0_230 (.A1(n_32_0_196), .A2(rst), .ZN(n_32_32));
   AOI22_X1 i_32_0_231 (.A1(n_32_0_4), .A2(\MEM[9] [17]), .B1(n_32_0_6), 
      .B2(\MEM[10] [17]), .ZN(n_32_0_197));
   AOI22_X1 i_32_0_232 (.A1(n_32_0_9), .A2(\MEM[5] [17]), .B1(n_32_0_12), 
      .B2(\MEM[3] [17]), .ZN(n_32_0_198));
   AOI22_X1 i_32_0_233 (.A1(\MEM[6] [17]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [17]), .ZN(n_32_0_199));
   AOI22_X1 i_32_0_234 (.A1(\MEM[8] [17]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [17]), .ZN(n_32_0_200));
   NAND4_X1 i_32_0_235 (.A1(n_32_0_197), .A2(n_32_0_198), .A3(n_32_0_199), 
      .A4(n_32_0_200), .ZN(n_32_0_201));
   AOI221_X1 i_32_0_236 (.A(n_32_0_201), .B1(\MEM[2] [17]), .B2(n_32_0_22), 
      .C1(\MEM[0] [17]), .C2(n_32_0_23), .ZN(n_32_0_202));
   AOI22_X1 i_32_0_237 (.A1(\MEM[4] [17]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [17]), .ZN(n_32_0_203));
   AOI22_X1 i_32_0_238 (.A1(\MEM[1] [17]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [17]), .ZN(n_32_0_204));
   AOI22_X1 i_32_0_239 (.A1(\MEM[12] [17]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [17]), .ZN(n_32_0_205));
   NAND4_X1 i_32_0_240 (.A1(n_32_0_202), .A2(n_32_0_203), .A3(n_32_0_204), 
      .A4(n_32_0_205), .ZN(MEM[17]));
   OAI22_X1 i_32_0_241 (.A1(MEM[17]), .A2(we1), .B1(data1[17]), .B2(n_32_0_35), 
      .ZN(n_32_0_206));
   NOR2_X1 i_32_0_242 (.A1(n_32_0_206), .A2(rst), .ZN(n_32_33));
   AOI22_X1 i_32_0_243 (.A1(n_32_0_4), .A2(\MEM[9] [18]), .B1(n_32_0_6), 
      .B2(\MEM[10] [18]), .ZN(n_32_0_207));
   AOI22_X1 i_32_0_244 (.A1(n_32_0_9), .A2(\MEM[5] [18]), .B1(n_32_0_12), 
      .B2(\MEM[3] [18]), .ZN(n_32_0_208));
   AOI22_X1 i_32_0_245 (.A1(\MEM[6] [18]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [18]), .ZN(n_32_0_209));
   AOI22_X1 i_32_0_246 (.A1(\MEM[8] [18]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [18]), .ZN(n_32_0_210));
   NAND4_X1 i_32_0_247 (.A1(n_32_0_207), .A2(n_32_0_208), .A3(n_32_0_209), 
      .A4(n_32_0_210), .ZN(n_32_0_211));
   AOI221_X1 i_32_0_248 (.A(n_32_0_211), .B1(\MEM[2] [18]), .B2(n_32_0_22), 
      .C1(\MEM[0] [18]), .C2(n_32_0_23), .ZN(n_32_0_212));
   AOI22_X1 i_32_0_249 (.A1(\MEM[4] [18]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [18]), .ZN(n_32_0_213));
   AOI22_X1 i_32_0_250 (.A1(\MEM[1] [18]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [18]), .ZN(n_32_0_214));
   AOI22_X1 i_32_0_251 (.A1(\MEM[12] [18]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [18]), .ZN(n_32_0_215));
   NAND4_X1 i_32_0_252 (.A1(n_32_0_212), .A2(n_32_0_213), .A3(n_32_0_214), 
      .A4(n_32_0_215), .ZN(MEM[18]));
   OAI22_X1 i_32_0_253 (.A1(MEM[18]), .A2(we1), .B1(data1[18]), .B2(n_32_0_35), 
      .ZN(n_32_0_216));
   NOR2_X1 i_32_0_254 (.A1(n_32_0_216), .A2(rst), .ZN(n_32_34));
   AOI22_X1 i_32_0_255 (.A1(n_32_0_4), .A2(\MEM[9] [19]), .B1(n_32_0_6), 
      .B2(\MEM[10] [19]), .ZN(n_32_0_217));
   AOI22_X1 i_32_0_256 (.A1(n_32_0_9), .A2(\MEM[5] [19]), .B1(n_32_0_12), 
      .B2(\MEM[3] [19]), .ZN(n_32_0_218));
   AOI22_X1 i_32_0_257 (.A1(\MEM[6] [19]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [19]), .ZN(n_32_0_219));
   AOI22_X1 i_32_0_258 (.A1(\MEM[8] [19]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [19]), .ZN(n_32_0_220));
   NAND4_X1 i_32_0_259 (.A1(n_32_0_217), .A2(n_32_0_218), .A3(n_32_0_219), 
      .A4(n_32_0_220), .ZN(n_32_0_221));
   AOI221_X1 i_32_0_260 (.A(n_32_0_221), .B1(\MEM[2] [19]), .B2(n_32_0_22), 
      .C1(\MEM[0] [19]), .C2(n_32_0_23), .ZN(n_32_0_222));
   AOI22_X1 i_32_0_261 (.A1(\MEM[4] [19]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [19]), .ZN(n_32_0_223));
   AOI22_X1 i_32_0_262 (.A1(\MEM[1] [19]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [19]), .ZN(n_32_0_224));
   AOI22_X1 i_32_0_263 (.A1(\MEM[12] [19]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [19]), .ZN(n_32_0_225));
   NAND4_X1 i_32_0_264 (.A1(n_32_0_222), .A2(n_32_0_223), .A3(n_32_0_224), 
      .A4(n_32_0_225), .ZN(MEM[19]));
   OAI22_X1 i_32_0_265 (.A1(MEM[19]), .A2(we1), .B1(data1[19]), .B2(n_32_0_35), 
      .ZN(n_32_0_226));
   NOR2_X1 i_32_0_266 (.A1(n_32_0_226), .A2(rst), .ZN(n_32_35));
   AOI22_X1 i_32_0_267 (.A1(n_32_0_4), .A2(\MEM[9] [20]), .B1(n_32_0_6), 
      .B2(\MEM[10] [20]), .ZN(n_32_0_227));
   AOI22_X1 i_32_0_268 (.A1(n_32_0_9), .A2(\MEM[5] [20]), .B1(n_32_0_12), 
      .B2(\MEM[3] [20]), .ZN(n_32_0_228));
   AOI22_X1 i_32_0_269 (.A1(\MEM[6] [20]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [20]), .ZN(n_32_0_229));
   AOI22_X1 i_32_0_270 (.A1(\MEM[8] [20]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [20]), .ZN(n_32_0_230));
   NAND4_X1 i_32_0_271 (.A1(n_32_0_227), .A2(n_32_0_228), .A3(n_32_0_229), 
      .A4(n_32_0_230), .ZN(n_32_0_231));
   AOI221_X1 i_32_0_272 (.A(n_32_0_231), .B1(\MEM[2] [20]), .B2(n_32_0_22), 
      .C1(\MEM[0] [20]), .C2(n_32_0_23), .ZN(n_32_0_232));
   AOI22_X1 i_32_0_273 (.A1(\MEM[4] [20]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [20]), .ZN(n_32_0_233));
   AOI22_X1 i_32_0_274 (.A1(\MEM[1] [20]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [20]), .ZN(n_32_0_234));
   AOI22_X1 i_32_0_275 (.A1(\MEM[12] [20]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [20]), .ZN(n_32_0_235));
   NAND4_X1 i_32_0_276 (.A1(n_32_0_232), .A2(n_32_0_233), .A3(n_32_0_234), 
      .A4(n_32_0_235), .ZN(MEM[20]));
   OAI22_X1 i_32_0_277 (.A1(MEM[20]), .A2(we1), .B1(data1[20]), .B2(n_32_0_35), 
      .ZN(n_32_0_236));
   NOR2_X1 i_32_0_278 (.A1(n_32_0_236), .A2(rst), .ZN(n_32_36));
   AOI22_X1 i_32_0_279 (.A1(n_32_0_4), .A2(\MEM[9] [21]), .B1(n_32_0_6), 
      .B2(\MEM[10] [21]), .ZN(n_32_0_237));
   AOI22_X1 i_32_0_280 (.A1(n_32_0_9), .A2(\MEM[5] [21]), .B1(n_32_0_12), 
      .B2(\MEM[3] [21]), .ZN(n_32_0_238));
   AOI22_X1 i_32_0_281 (.A1(\MEM[6] [21]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [21]), .ZN(n_32_0_239));
   AOI22_X1 i_32_0_282 (.A1(\MEM[8] [21]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [21]), .ZN(n_32_0_240));
   NAND4_X1 i_32_0_283 (.A1(n_32_0_237), .A2(n_32_0_238), .A3(n_32_0_239), 
      .A4(n_32_0_240), .ZN(n_32_0_241));
   AOI221_X1 i_32_0_284 (.A(n_32_0_241), .B1(\MEM[2] [21]), .B2(n_32_0_22), 
      .C1(\MEM[0] [21]), .C2(n_32_0_23), .ZN(n_32_0_242));
   AOI22_X1 i_32_0_285 (.A1(\MEM[4] [21]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [21]), .ZN(n_32_0_243));
   AOI22_X1 i_32_0_286 (.A1(\MEM[1] [21]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [21]), .ZN(n_32_0_244));
   AOI22_X1 i_32_0_287 (.A1(\MEM[12] [21]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [21]), .ZN(n_32_0_245));
   NAND4_X1 i_32_0_288 (.A1(n_32_0_242), .A2(n_32_0_243), .A3(n_32_0_244), 
      .A4(n_32_0_245), .ZN(MEM[21]));
   OAI22_X1 i_32_0_289 (.A1(MEM[21]), .A2(we1), .B1(data1[21]), .B2(n_32_0_35), 
      .ZN(n_32_0_246));
   NOR2_X1 i_32_0_290 (.A1(n_32_0_246), .A2(rst), .ZN(n_32_37));
   AOI22_X1 i_32_0_291 (.A1(n_32_0_4), .A2(\MEM[9] [22]), .B1(n_32_0_6), 
      .B2(\MEM[10] [22]), .ZN(n_32_0_247));
   AOI22_X1 i_32_0_292 (.A1(n_32_0_9), .A2(\MEM[5] [22]), .B1(n_32_0_12), 
      .B2(\MEM[3] [22]), .ZN(n_32_0_248));
   AOI22_X1 i_32_0_293 (.A1(\MEM[6] [22]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [22]), .ZN(n_32_0_249));
   AOI22_X1 i_32_0_294 (.A1(\MEM[8] [22]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [22]), .ZN(n_32_0_250));
   NAND4_X1 i_32_0_295 (.A1(n_32_0_247), .A2(n_32_0_248), .A3(n_32_0_249), 
      .A4(n_32_0_250), .ZN(n_32_0_251));
   AOI221_X1 i_32_0_296 (.A(n_32_0_251), .B1(\MEM[2] [22]), .B2(n_32_0_22), 
      .C1(\MEM[0] [22]), .C2(n_32_0_23), .ZN(n_32_0_252));
   AOI22_X1 i_32_0_297 (.A1(\MEM[4] [22]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [22]), .ZN(n_32_0_253));
   AOI22_X1 i_32_0_298 (.A1(\MEM[1] [22]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [22]), .ZN(n_32_0_254));
   AOI22_X1 i_32_0_299 (.A1(\MEM[12] [22]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [22]), .ZN(n_32_0_255));
   NAND4_X1 i_32_0_300 (.A1(n_32_0_252), .A2(n_32_0_253), .A3(n_32_0_254), 
      .A4(n_32_0_255), .ZN(MEM[22]));
   OAI22_X1 i_32_0_301 (.A1(MEM[22]), .A2(we1), .B1(data1[22]), .B2(n_32_0_35), 
      .ZN(n_32_0_256));
   NOR2_X1 i_32_0_302 (.A1(n_32_0_256), .A2(rst), .ZN(n_32_38));
   AOI22_X1 i_32_0_303 (.A1(n_32_0_4), .A2(\MEM[9] [23]), .B1(n_32_0_6), 
      .B2(\MEM[10] [23]), .ZN(n_32_0_257));
   AOI22_X1 i_32_0_304 (.A1(n_32_0_9), .A2(\MEM[5] [23]), .B1(n_32_0_12), 
      .B2(\MEM[3] [23]), .ZN(n_32_0_258));
   AOI22_X1 i_32_0_305 (.A1(\MEM[6] [23]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [23]), .ZN(n_32_0_259));
   AOI22_X1 i_32_0_306 (.A1(\MEM[8] [23]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [23]), .ZN(n_32_0_260));
   NAND4_X1 i_32_0_307 (.A1(n_32_0_257), .A2(n_32_0_258), .A3(n_32_0_259), 
      .A4(n_32_0_260), .ZN(n_32_0_261));
   AOI221_X1 i_32_0_308 (.A(n_32_0_261), .B1(\MEM[2] [23]), .B2(n_32_0_22), 
      .C1(\MEM[0] [23]), .C2(n_32_0_23), .ZN(n_32_0_262));
   AOI22_X1 i_32_0_309 (.A1(\MEM[4] [23]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [23]), .ZN(n_32_0_263));
   AOI22_X1 i_32_0_310 (.A1(\MEM[1] [23]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [23]), .ZN(n_32_0_264));
   AOI22_X1 i_32_0_311 (.A1(\MEM[12] [23]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [23]), .ZN(n_32_0_265));
   NAND4_X1 i_32_0_312 (.A1(n_32_0_262), .A2(n_32_0_263), .A3(n_32_0_264), 
      .A4(n_32_0_265), .ZN(MEM[23]));
   OAI22_X1 i_32_0_313 (.A1(MEM[23]), .A2(we1), .B1(data1[23]), .B2(n_32_0_35), 
      .ZN(n_32_0_266));
   NOR2_X1 i_32_0_314 (.A1(n_32_0_266), .A2(rst), .ZN(n_32_39));
   AOI22_X1 i_32_0_315 (.A1(n_32_0_4), .A2(\MEM[9] [24]), .B1(n_32_0_6), 
      .B2(\MEM[10] [24]), .ZN(n_32_0_267));
   AOI22_X1 i_32_0_316 (.A1(n_32_0_9), .A2(\MEM[5] [24]), .B1(n_32_0_12), 
      .B2(\MEM[3] [24]), .ZN(n_32_0_268));
   AOI22_X1 i_32_0_317 (.A1(\MEM[6] [24]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [24]), .ZN(n_32_0_269));
   AOI22_X1 i_32_0_318 (.A1(\MEM[8] [24]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [24]), .ZN(n_32_0_270));
   NAND4_X1 i_32_0_319 (.A1(n_32_0_267), .A2(n_32_0_268), .A3(n_32_0_269), 
      .A4(n_32_0_270), .ZN(n_32_0_271));
   AOI221_X1 i_32_0_320 (.A(n_32_0_271), .B1(\MEM[2] [24]), .B2(n_32_0_22), 
      .C1(\MEM[0] [24]), .C2(n_32_0_23), .ZN(n_32_0_272));
   AOI22_X1 i_32_0_321 (.A1(\MEM[4] [24]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [24]), .ZN(n_32_0_273));
   AOI22_X1 i_32_0_322 (.A1(\MEM[1] [24]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [24]), .ZN(n_32_0_274));
   AOI22_X1 i_32_0_323 (.A1(\MEM[12] [24]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [24]), .ZN(n_32_0_275));
   NAND4_X1 i_32_0_324 (.A1(n_32_0_272), .A2(n_32_0_273), .A3(n_32_0_274), 
      .A4(n_32_0_275), .ZN(MEM[24]));
   OAI22_X1 i_32_0_325 (.A1(MEM[24]), .A2(we1), .B1(data1[24]), .B2(n_32_0_35), 
      .ZN(n_32_0_276));
   NOR2_X1 i_32_0_326 (.A1(n_32_0_276), .A2(rst), .ZN(n_32_40));
   AOI22_X1 i_32_0_327 (.A1(n_32_0_4), .A2(\MEM[9] [25]), .B1(n_32_0_6), 
      .B2(\MEM[10] [25]), .ZN(n_32_0_277));
   AOI22_X1 i_32_0_328 (.A1(n_32_0_9), .A2(\MEM[5] [25]), .B1(n_32_0_12), 
      .B2(\MEM[3] [25]), .ZN(n_32_0_278));
   AOI22_X1 i_32_0_329 (.A1(\MEM[6] [25]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [25]), .ZN(n_32_0_279));
   AOI22_X1 i_32_0_330 (.A1(\MEM[8] [25]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [25]), .ZN(n_32_0_280));
   NAND4_X1 i_32_0_331 (.A1(n_32_0_277), .A2(n_32_0_278), .A3(n_32_0_279), 
      .A4(n_32_0_280), .ZN(n_32_0_281));
   AOI221_X1 i_32_0_332 (.A(n_32_0_281), .B1(\MEM[2] [25]), .B2(n_32_0_22), 
      .C1(\MEM[0] [25]), .C2(n_32_0_23), .ZN(n_32_0_282));
   AOI22_X1 i_32_0_333 (.A1(\MEM[4] [25]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [25]), .ZN(n_32_0_283));
   AOI22_X1 i_32_0_334 (.A1(\MEM[1] [25]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [25]), .ZN(n_32_0_284));
   AOI22_X1 i_32_0_335 (.A1(\MEM[12] [25]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [25]), .ZN(n_32_0_285));
   NAND4_X1 i_32_0_336 (.A1(n_32_0_282), .A2(n_32_0_283), .A3(n_32_0_284), 
      .A4(n_32_0_285), .ZN(MEM[25]));
   OAI22_X1 i_32_0_337 (.A1(MEM[25]), .A2(we1), .B1(data1[25]), .B2(n_32_0_35), 
      .ZN(n_32_0_286));
   NOR2_X1 i_32_0_338 (.A1(n_32_0_286), .A2(rst), .ZN(n_32_41));
   AOI22_X1 i_32_0_339 (.A1(n_32_0_4), .A2(\MEM[9] [26]), .B1(n_32_0_6), 
      .B2(\MEM[10] [26]), .ZN(n_32_0_287));
   AOI22_X1 i_32_0_340 (.A1(n_32_0_9), .A2(\MEM[5] [26]), .B1(n_32_0_12), 
      .B2(\MEM[3] [26]), .ZN(n_32_0_288));
   AOI22_X1 i_32_0_341 (.A1(\MEM[6] [26]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [26]), .ZN(n_32_0_289));
   AOI22_X1 i_32_0_342 (.A1(\MEM[8] [26]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [26]), .ZN(n_32_0_290));
   NAND4_X1 i_32_0_343 (.A1(n_32_0_287), .A2(n_32_0_288), .A3(n_32_0_289), 
      .A4(n_32_0_290), .ZN(n_32_0_291));
   AOI221_X1 i_32_0_344 (.A(n_32_0_291), .B1(\MEM[2] [26]), .B2(n_32_0_22), 
      .C1(\MEM[0] [26]), .C2(n_32_0_23), .ZN(n_32_0_292));
   AOI22_X1 i_32_0_345 (.A1(\MEM[4] [26]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [26]), .ZN(n_32_0_293));
   AOI22_X1 i_32_0_346 (.A1(\MEM[1] [26]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [26]), .ZN(n_32_0_294));
   AOI22_X1 i_32_0_347 (.A1(\MEM[12] [26]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [26]), .ZN(n_32_0_295));
   NAND4_X1 i_32_0_348 (.A1(n_32_0_292), .A2(n_32_0_293), .A3(n_32_0_294), 
      .A4(n_32_0_295), .ZN(MEM[26]));
   OAI22_X1 i_32_0_349 (.A1(MEM[26]), .A2(we1), .B1(data1[26]), .B2(n_32_0_35), 
      .ZN(n_32_0_296));
   NOR2_X1 i_32_0_350 (.A1(n_32_0_296), .A2(rst), .ZN(n_32_42));
   AOI22_X1 i_32_0_351 (.A1(n_32_0_4), .A2(\MEM[9] [27]), .B1(n_32_0_6), 
      .B2(\MEM[10] [27]), .ZN(n_32_0_297));
   AOI22_X1 i_32_0_352 (.A1(n_32_0_9), .A2(\MEM[5] [27]), .B1(n_32_0_12), 
      .B2(\MEM[3] [27]), .ZN(n_32_0_298));
   AOI22_X1 i_32_0_353 (.A1(\MEM[6] [27]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [27]), .ZN(n_32_0_299));
   AOI22_X1 i_32_0_354 (.A1(\MEM[8] [27]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [27]), .ZN(n_32_0_300));
   NAND4_X1 i_32_0_355 (.A1(n_32_0_297), .A2(n_32_0_298), .A3(n_32_0_299), 
      .A4(n_32_0_300), .ZN(n_32_0_301));
   AOI221_X1 i_32_0_356 (.A(n_32_0_301), .B1(\MEM[2] [27]), .B2(n_32_0_22), 
      .C1(\MEM[0] [27]), .C2(n_32_0_23), .ZN(n_32_0_302));
   AOI22_X1 i_32_0_357 (.A1(\MEM[4] [27]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [27]), .ZN(n_32_0_303));
   AOI22_X1 i_32_0_358 (.A1(\MEM[1] [27]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [27]), .ZN(n_32_0_304));
   AOI22_X1 i_32_0_359 (.A1(\MEM[12] [27]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [27]), .ZN(n_32_0_305));
   NAND4_X1 i_32_0_360 (.A1(n_32_0_302), .A2(n_32_0_303), .A3(n_32_0_304), 
      .A4(n_32_0_305), .ZN(MEM[27]));
   OAI22_X1 i_32_0_361 (.A1(MEM[27]), .A2(we1), .B1(data1[27]), .B2(n_32_0_35), 
      .ZN(n_32_0_306));
   NOR2_X1 i_32_0_362 (.A1(n_32_0_306), .A2(rst), .ZN(n_32_43));
   AOI22_X1 i_32_0_363 (.A1(n_32_0_4), .A2(\MEM[9] [28]), .B1(n_32_0_6), 
      .B2(\MEM[10] [28]), .ZN(n_32_0_307));
   AOI22_X1 i_32_0_364 (.A1(n_32_0_9), .A2(\MEM[5] [28]), .B1(n_32_0_12), 
      .B2(\MEM[3] [28]), .ZN(n_32_0_308));
   AOI22_X1 i_32_0_365 (.A1(\MEM[6] [28]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [28]), .ZN(n_32_0_309));
   AOI22_X1 i_32_0_366 (.A1(\MEM[8] [28]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [28]), .ZN(n_32_0_310));
   NAND4_X1 i_32_0_367 (.A1(n_32_0_307), .A2(n_32_0_308), .A3(n_32_0_309), 
      .A4(n_32_0_310), .ZN(n_32_0_311));
   AOI221_X1 i_32_0_368 (.A(n_32_0_311), .B1(\MEM[2] [28]), .B2(n_32_0_22), 
      .C1(\MEM[0] [28]), .C2(n_32_0_23), .ZN(n_32_0_312));
   AOI22_X1 i_32_0_369 (.A1(\MEM[4] [28]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [28]), .ZN(n_32_0_313));
   AOI22_X1 i_32_0_370 (.A1(\MEM[1] [28]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [28]), .ZN(n_32_0_314));
   AOI22_X1 i_32_0_371 (.A1(\MEM[12] [28]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [28]), .ZN(n_32_0_315));
   NAND4_X1 i_32_0_372 (.A1(n_32_0_312), .A2(n_32_0_313), .A3(n_32_0_314), 
      .A4(n_32_0_315), .ZN(MEM[28]));
   OAI22_X1 i_32_0_373 (.A1(MEM[28]), .A2(we1), .B1(data1[28]), .B2(n_32_0_35), 
      .ZN(n_32_0_316));
   NOR2_X1 i_32_0_374 (.A1(n_32_0_316), .A2(rst), .ZN(n_32_44));
   AOI22_X1 i_32_0_375 (.A1(n_32_0_4), .A2(\MEM[9] [29]), .B1(n_32_0_6), 
      .B2(\MEM[10] [29]), .ZN(n_32_0_317));
   AOI22_X1 i_32_0_376 (.A1(n_32_0_9), .A2(\MEM[5] [29]), .B1(n_32_0_12), 
      .B2(\MEM[3] [29]), .ZN(n_32_0_318));
   AOI22_X1 i_32_0_377 (.A1(\MEM[6] [29]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [29]), .ZN(n_32_0_319));
   AOI22_X1 i_32_0_378 (.A1(\MEM[8] [29]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [29]), .ZN(n_32_0_320));
   NAND4_X1 i_32_0_379 (.A1(n_32_0_317), .A2(n_32_0_318), .A3(n_32_0_319), 
      .A4(n_32_0_320), .ZN(n_32_0_321));
   AOI221_X1 i_32_0_380 (.A(n_32_0_321), .B1(\MEM[2] [29]), .B2(n_32_0_22), 
      .C1(\MEM[0] [29]), .C2(n_32_0_23), .ZN(n_32_0_322));
   AOI22_X1 i_32_0_381 (.A1(\MEM[4] [29]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [29]), .ZN(n_32_0_323));
   AOI22_X1 i_32_0_382 (.A1(\MEM[1] [29]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [29]), .ZN(n_32_0_324));
   AOI22_X1 i_32_0_383 (.A1(\MEM[12] [29]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [29]), .ZN(n_32_0_325));
   NAND4_X1 i_32_0_384 (.A1(n_32_0_322), .A2(n_32_0_323), .A3(n_32_0_324), 
      .A4(n_32_0_325), .ZN(MEM[29]));
   OAI22_X1 i_32_0_385 (.A1(MEM[29]), .A2(we1), .B1(data1[29]), .B2(n_32_0_35), 
      .ZN(n_32_0_326));
   NOR2_X1 i_32_0_386 (.A1(n_32_0_326), .A2(rst), .ZN(n_32_45));
   AOI22_X1 i_32_0_387 (.A1(n_32_0_4), .A2(\MEM[9] [30]), .B1(n_32_0_6), 
      .B2(\MEM[10] [30]), .ZN(n_32_0_327));
   AOI22_X1 i_32_0_388 (.A1(n_32_0_9), .A2(\MEM[5] [30]), .B1(n_32_0_12), 
      .B2(\MEM[3] [30]), .ZN(n_32_0_328));
   AOI22_X1 i_32_0_389 (.A1(\MEM[6] [30]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [30]), .ZN(n_32_0_329));
   AOI22_X1 i_32_0_390 (.A1(\MEM[8] [30]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [30]), .ZN(n_32_0_330));
   NAND4_X1 i_32_0_391 (.A1(n_32_0_327), .A2(n_32_0_328), .A3(n_32_0_329), 
      .A4(n_32_0_330), .ZN(n_32_0_331));
   AOI221_X1 i_32_0_392 (.A(n_32_0_331), .B1(\MEM[2] [30]), .B2(n_32_0_22), 
      .C1(\MEM[0] [30]), .C2(n_32_0_23), .ZN(n_32_0_332));
   AOI22_X1 i_32_0_393 (.A1(\MEM[4] [30]), .A2(n_32_0_25), .B1(n_32_0_27), 
      .B2(\MEM[13] [30]), .ZN(n_32_0_333));
   AOI22_X1 i_32_0_394 (.A1(\MEM[1] [30]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [30]), .ZN(n_32_0_334));
   AOI22_X1 i_32_0_395 (.A1(\MEM[12] [30]), .A2(n_32_0_32), .B1(n_32_0_33), 
      .B2(\MEM[14] [30]), .ZN(n_32_0_335));
   NAND4_X1 i_32_0_396 (.A1(n_32_0_332), .A2(n_32_0_333), .A3(n_32_0_334), 
      .A4(n_32_0_335), .ZN(MEM[30]));
   OAI22_X1 i_32_0_397 (.A1(MEM[30]), .A2(we1), .B1(data1[30]), .B2(n_32_0_35), 
      .ZN(n_32_0_336));
   NOR2_X1 i_32_0_398 (.A1(n_32_0_336), .A2(rst), .ZN(n_32_46));
   INV_X1 i_32_0_399 (.A(data1[31]), .ZN(n_32_0_337));
   AOI22_X1 i_32_0_400 (.A1(\MEM[2] [31]), .A2(n_32_0_22), .B1(n_32_0_9), 
      .B2(\MEM[5] [31]), .ZN(n_32_0_338));
   AOI22_X1 i_32_0_401 (.A1(n_32_0_6), .A2(\MEM[10] [31]), .B1(n_32_0_4), 
      .B2(\MEM[9] [31]), .ZN(n_32_0_339));
   AOI22_X1 i_32_0_402 (.A1(\MEM[4] [31]), .A2(n_32_0_25), .B1(n_32_0_12), 
      .B2(\MEM[3] [31]), .ZN(n_32_0_340));
   AOI22_X1 i_32_0_403 (.A1(n_32_0_23), .A2(\MEM[0] [31]), .B1(n_32_0_33), 
      .B2(\MEM[14] [31]), .ZN(n_32_0_341));
   NAND4_X1 i_32_0_404 (.A1(n_32_0_338), .A2(n_32_0_339), .A3(n_32_0_340), 
      .A4(n_32_0_341), .ZN(n_32_0_342));
   AOI22_X1 i_32_0_405 (.A1(n_32_0_32), .A2(\MEM[12] [31]), .B1(n_32_0_27), 
      .B2(\MEM[13] [31]), .ZN(n_32_0_343));
   AOI22_X1 i_32_0_406 (.A1(\MEM[8] [31]), .A2(n_32_0_18), .B1(n_32_0_19), 
      .B2(\MEM[11] [31]), .ZN(n_32_0_344));
   AOI22_X1 i_32_0_407 (.A1(\MEM[6] [31]), .A2(n_32_0_14), .B1(n_32_0_15), 
      .B2(\MEM[7] [31]), .ZN(n_32_0_345));
   AOI22_X1 i_32_0_408 (.A1(\MEM[1] [31]), .A2(n_32_0_29), .B1(n_32_0_30), 
      .B2(\MEM[15] [31]), .ZN(n_32_0_346));
   NAND4_X1 i_32_0_409 (.A1(n_32_0_343), .A2(n_32_0_344), .A3(n_32_0_345), 
      .A4(n_32_0_346), .ZN(n_32_0_347));
   NOR2_X1 i_32_0_410 (.A1(n_32_0_342), .A2(n_32_0_347), .ZN(n_32_0_348));
   AOI221_X1 i_32_0_411 (.A(rst), .B1(n_32_0_337), .B2(we1), .C1(n_32_0_348), 
      .C2(n_32_0_35), .ZN(n_32_47));
   OR2_X1 i_32_0_412 (.A1(n_32_0_23), .A2(rst), .ZN(n_32_48));
   OR2_X1 i_32_0_413 (.A1(n_32_0_29), .A2(rst), .ZN(n_32_49));
   OR2_X1 i_32_0_414 (.A1(n_32_0_22), .A2(rst), .ZN(n_32_50));
   OR2_X1 i_32_0_415 (.A1(n_32_0_12), .A2(rst), .ZN(n_32_51));
   OR2_X1 i_32_0_416 (.A1(n_32_0_25), .A2(rst), .ZN(n_32_52));
   OR2_X1 i_32_0_417 (.A1(n_32_0_9), .A2(rst), .ZN(n_32_53));
   OR2_X1 i_32_0_418 (.A1(n_32_0_14), .A2(rst), .ZN(n_32_54));
   OR2_X1 i_32_0_419 (.A1(n_32_0_15), .A2(rst), .ZN(n_32_55));
   OR2_X1 i_32_0_420 (.A1(n_32_0_18), .A2(rst), .ZN(n_32_56));
   OR2_X1 i_32_0_421 (.A1(n_32_0_4), .A2(rst), .ZN(n_32_57));
   OR2_X1 i_32_0_422 (.A1(n_32_0_6), .A2(rst), .ZN(n_32_58));
   OR2_X1 i_32_0_423 (.A1(n_32_0_19), .A2(rst), .ZN(n_32_59));
   OR2_X1 i_32_0_424 (.A1(n_32_0_32), .A2(rst), .ZN(n_32_60));
   OR2_X1 i_32_0_425 (.A1(n_32_0_27), .A2(rst), .ZN(n_32_61));
   OR2_X1 i_32_0_426 (.A1(n_32_0_33), .A2(rst), .ZN(n_32_62));
   OR2_X1 i_32_0_427 (.A1(n_32_0_30), .A2(rst), .ZN(n_32_63));
   INV_X1 i_32_0_428 (.A(addr2[0]), .ZN(n_32_0_349));
   INV_X1 i_32_0_429 (.A(addr2[1]), .ZN(n_32_0_350));
   NAND2_X1 i_32_0_430 (.A1(n_32_0_349), .A2(n_32_0_350), .ZN(n_32_0_351));
   INV_X1 i_32_0_431 (.A(addr2[3]), .ZN(n_32_0_352));
   INV_X1 i_32_0_432 (.A(addr2[2]), .ZN(n_32_0_353));
   NAND2_X1 i_32_0_433 (.A1(n_32_0_352), .A2(n_32_0_353), .ZN(n_32_0_354));
   NOR2_X1 i_32_0_434 (.A1(n_32_0_351), .A2(n_32_0_354), .ZN(n_32_0_355));
   NAND2_X1 i_32_0_435 (.A1(n_32_0_349), .A2(addr2[1]), .ZN(n_32_0_356));
   NOR2_X1 i_32_0_436 (.A1(n_32_0_354), .A2(n_32_0_356), .ZN(n_32_0_357));
   AOI22_X1 i_32_0_437 (.A1(n_32_0_355), .A2(\MEM[0] [0]), .B1(n_32_0_357), 
      .B2(\MEM[2] [0]), .ZN(n_32_0_358));
   NAND2_X1 i_32_0_438 (.A1(n_32_0_352), .A2(addr2[2]), .ZN(n_32_0_359));
   NOR2_X1 i_32_0_439 (.A1(n_32_0_351), .A2(n_32_0_359), .ZN(n_32_0_360));
   NAND2_X1 i_32_0_440 (.A1(n_32_0_350), .A2(addr2[0]), .ZN(n_32_0_361));
   NAND2_X1 i_32_0_441 (.A1(addr2[3]), .A2(addr2[2]), .ZN(n_32_0_362));
   NOR2_X1 i_32_0_442 (.A1(n_32_0_361), .A2(n_32_0_362), .ZN(n_32_0_363));
   AOI22_X1 i_32_0_443 (.A1(\MEM[4] [0]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [0]), .ZN(n_32_0_364));
   NOR2_X1 i_32_0_444 (.A1(n_32_0_351), .A2(n_32_0_362), .ZN(n_32_0_365));
   NOR2_X1 i_32_0_445 (.A1(n_32_0_356), .A2(n_32_0_362), .ZN(n_32_0_366));
   AOI22_X1 i_32_0_446 (.A1(\MEM[12] [0]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [0]), .ZN(n_32_0_367));
   NOR2_X1 i_32_0_447 (.A1(n_32_0_354), .A2(n_32_0_361), .ZN(n_32_0_368));
   NAND2_X1 i_32_0_448 (.A1(addr2[0]), .A2(addr2[1]), .ZN(n_32_0_369));
   NOR2_X1 i_32_0_449 (.A1(n_32_0_369), .A2(n_32_0_362), .ZN(n_32_0_370));
   AOI22_X1 i_32_0_450 (.A1(\MEM[1] [0]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [0]), .ZN(n_32_0_371));
   NAND4_X1 i_32_0_451 (.A1(n_32_0_358), .A2(n_32_0_364), .A3(n_32_0_367), 
      .A4(n_32_0_371), .ZN(n_32_0_372));
   NAND2_X1 i_32_0_452 (.A1(n_32_0_353), .A2(addr2[3]), .ZN(n_32_0_373));
   NOR2_X1 i_32_0_453 (.A1(n_32_0_373), .A2(n_32_0_361), .ZN(n_32_0_374));
   NOR2_X1 i_32_0_454 (.A1(n_32_0_373), .A2(n_32_0_356), .ZN(n_32_0_375));
   AOI221_X1 i_32_0_455 (.A(n_32_0_372), .B1(\MEM[9] [0]), .B2(n_32_0_374), 
      .C1(\MEM[10] [0]), .C2(n_32_0_375), .ZN(n_32_0_376));
   NOR2_X1 i_32_0_456 (.A1(n_32_0_351), .A2(n_32_0_373), .ZN(n_32_0_377));
   NOR2_X1 i_32_0_457 (.A1(n_32_0_373), .A2(n_32_0_369), .ZN(n_32_0_378));
   AOI22_X1 i_32_0_458 (.A1(\MEM[8] [0]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [0]), .ZN(n_32_0_379));
   NOR2_X1 i_32_0_459 (.A1(n_32_0_359), .A2(n_32_0_356), .ZN(n_32_0_380));
   NOR2_X1 i_32_0_460 (.A1(n_32_0_359), .A2(n_32_0_369), .ZN(n_32_0_381));
   AOI22_X1 i_32_0_461 (.A1(\MEM[6] [0]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [0]), .ZN(n_32_0_382));
   NOR2_X1 i_32_0_462 (.A1(n_32_0_359), .A2(n_32_0_361), .ZN(n_32_0_383));
   NOR2_X1 i_32_0_463 (.A1(n_32_0_354), .A2(n_32_0_369), .ZN(n_32_0_384));
   AOI22_X1 i_32_0_464 (.A1(n_32_0_383), .A2(\MEM[5] [0]), .B1(n_32_0_384), 
      .B2(\MEM[3] [0]), .ZN(n_32_0_385));
   NAND4_X1 i_32_0_465 (.A1(n_32_0_376), .A2(n_32_0_379), .A3(n_32_0_382), 
      .A4(n_32_0_385), .ZN(data2[0]));
   AOI22_X1 i_32_0_466 (.A1(n_32_0_355), .A2(\MEM[0] [1]), .B1(n_32_0_357), 
      .B2(\MEM[2] [1]), .ZN(n_32_0_386));
   AOI22_X1 i_32_0_467 (.A1(\MEM[4] [1]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [1]), .ZN(n_32_0_387));
   AOI22_X1 i_32_0_468 (.A1(n_32_0_365), .A2(\MEM[12] [1]), .B1(n_32_0_366), 
      .B2(\MEM[14] [1]), .ZN(n_32_0_388));
   AOI22_X1 i_32_0_469 (.A1(n_32_0_368), .A2(\MEM[1] [1]), .B1(n_32_0_370), 
      .B2(\MEM[15] [1]), .ZN(n_32_0_389));
   NAND4_X1 i_32_0_470 (.A1(n_32_0_386), .A2(n_32_0_387), .A3(n_32_0_388), 
      .A4(n_32_0_389), .ZN(n_32_0_390));
   AOI221_X1 i_32_0_471 (.A(n_32_0_390), .B1(\MEM[9] [1]), .B2(n_32_0_374), 
      .C1(\MEM[10] [1]), .C2(n_32_0_375), .ZN(n_32_0_391));
   AOI22_X1 i_32_0_472 (.A1(\MEM[8] [1]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [1]), .ZN(n_32_0_392));
   AOI22_X1 i_32_0_473 (.A1(\MEM[5] [1]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [1]), .ZN(n_32_0_393));
   AOI22_X1 i_32_0_474 (.A1(\MEM[6] [1]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [1]), .ZN(n_32_0_394));
   NAND4_X1 i_32_0_475 (.A1(n_32_0_391), .A2(n_32_0_392), .A3(n_32_0_393), 
      .A4(n_32_0_394), .ZN(data2[1]));
   AOI22_X1 i_32_0_476 (.A1(n_32_0_355), .A2(\MEM[0] [2]), .B1(n_32_0_357), 
      .B2(\MEM[2] [2]), .ZN(n_32_0_395));
   AOI22_X1 i_32_0_477 (.A1(n_32_0_360), .A2(\MEM[4] [2]), .B1(n_32_0_363), 
      .B2(\MEM[13] [2]), .ZN(n_32_0_396));
   AOI22_X1 i_32_0_478 (.A1(n_32_0_365), .A2(\MEM[12] [2]), .B1(n_32_0_366), 
      .B2(\MEM[14] [2]), .ZN(n_32_0_397));
   AOI22_X1 i_32_0_479 (.A1(n_32_0_368), .A2(\MEM[1] [2]), .B1(n_32_0_370), 
      .B2(\MEM[15] [2]), .ZN(n_32_0_398));
   NAND4_X1 i_32_0_480 (.A1(n_32_0_395), .A2(n_32_0_396), .A3(n_32_0_397), 
      .A4(n_32_0_398), .ZN(n_32_0_399));
   AOI221_X1 i_32_0_481 (.A(n_32_0_399), .B1(\MEM[10] [2]), .B2(n_32_0_375), 
      .C1(\MEM[9] [2]), .C2(n_32_0_374), .ZN(n_32_0_400));
   AOI22_X1 i_32_0_482 (.A1(n_32_0_380), .A2(\MEM[6] [2]), .B1(n_32_0_381), 
      .B2(\MEM[7] [2]), .ZN(n_32_0_401));
   AOI22_X1 i_32_0_483 (.A1(\MEM[8] [2]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [2]), .ZN(n_32_0_402));
   AOI22_X1 i_32_0_484 (.A1(\MEM[5] [2]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [2]), .ZN(n_32_0_403));
   NAND4_X1 i_32_0_485 (.A1(n_32_0_400), .A2(n_32_0_401), .A3(n_32_0_402), 
      .A4(n_32_0_403), .ZN(data2[2]));
   AOI22_X1 i_32_0_486 (.A1(\MEM[0] [3]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [3]), .ZN(n_32_0_404));
   AOI22_X1 i_32_0_487 (.A1(n_32_0_360), .A2(\MEM[4] [3]), .B1(n_32_0_363), 
      .B2(\MEM[13] [3]), .ZN(n_32_0_405));
   AOI22_X1 i_32_0_488 (.A1(\MEM[12] [3]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [3]), .ZN(n_32_0_406));
   AOI22_X1 i_32_0_489 (.A1(n_32_0_368), .A2(\MEM[1] [3]), .B1(n_32_0_370), 
      .B2(\MEM[15] [3]), .ZN(n_32_0_407));
   NAND4_X1 i_32_0_490 (.A1(n_32_0_404), .A2(n_32_0_405), .A3(n_32_0_406), 
      .A4(n_32_0_407), .ZN(n_32_0_408));
   AOI221_X1 i_32_0_491 (.A(n_32_0_408), .B1(\MEM[10] [3]), .B2(n_32_0_375), 
      .C1(\MEM[9] [3]), .C2(n_32_0_374), .ZN(n_32_0_409));
   AOI22_X1 i_32_0_492 (.A1(\MEM[8] [3]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [3]), .ZN(n_32_0_410));
   AOI22_X1 i_32_0_493 (.A1(n_32_0_380), .A2(\MEM[6] [3]), .B1(n_32_0_381), 
      .B2(\MEM[7] [3]), .ZN(n_32_0_411));
   AOI22_X1 i_32_0_494 (.A1(\MEM[5] [3]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [3]), .ZN(n_32_0_412));
   NAND4_X1 i_32_0_495 (.A1(n_32_0_409), .A2(n_32_0_410), .A3(n_32_0_411), 
      .A4(n_32_0_412), .ZN(data2[3]));
   AOI22_X1 i_32_0_496 (.A1(\MEM[0] [4]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [4]), .ZN(n_32_0_413));
   AOI22_X1 i_32_0_497 (.A1(n_32_0_360), .A2(\MEM[4] [4]), .B1(n_32_0_363), 
      .B2(\MEM[13] [4]), .ZN(n_32_0_414));
   NAND2_X1 i_32_0_498 (.A1(n_32_0_413), .A2(n_32_0_414), .ZN(n_32_0_415));
   AOI221_X1 i_32_0_499 (.A(n_32_0_415), .B1(\MEM[14] [4]), .B2(n_32_0_366), 
      .C1(\MEM[12] [4]), .C2(n_32_0_365), .ZN(n_32_0_416));
   AOI22_X1 i_32_0_500 (.A1(\MEM[5] [4]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [4]), .ZN(n_32_0_417));
   AOI22_X1 i_32_0_501 (.A1(n_32_0_380), .A2(\MEM[6] [4]), .B1(n_32_0_381), 
      .B2(\MEM[7] [4]), .ZN(n_32_0_418));
   NAND2_X1 i_32_0_502 (.A1(n_32_0_417), .A2(n_32_0_418), .ZN(n_32_0_419));
   AOI221_X1 i_32_0_503 (.A(n_32_0_419), .B1(\MEM[11] [4]), .B2(n_32_0_378), 
      .C1(\MEM[8] [4]), .C2(n_32_0_377), .ZN(n_32_0_420));
   AOI22_X1 i_32_0_504 (.A1(\MEM[1] [4]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [4]), .ZN(n_32_0_421));
   AOI22_X1 i_32_0_505 (.A1(n_32_0_375), .A2(\MEM[10] [4]), .B1(n_32_0_374), 
      .B2(\MEM[9] [4]), .ZN(n_32_0_422));
   NAND4_X1 i_32_0_506 (.A1(n_32_0_416), .A2(n_32_0_420), .A3(n_32_0_421), 
      .A4(n_32_0_422), .ZN(data2[4]));
   AOI22_X1 i_32_0_507 (.A1(n_32_0_355), .A2(\MEM[0] [5]), .B1(n_32_0_357), 
      .B2(\MEM[2] [5]), .ZN(n_32_0_423));
   AOI22_X1 i_32_0_508 (.A1(\MEM[4] [5]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [5]), .ZN(n_32_0_424));
   AOI22_X1 i_32_0_509 (.A1(\MEM[12] [5]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [5]), .ZN(n_32_0_425));
   AOI22_X1 i_32_0_510 (.A1(\MEM[1] [5]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [5]), .ZN(n_32_0_426));
   NAND4_X1 i_32_0_511 (.A1(n_32_0_423), .A2(n_32_0_424), .A3(n_32_0_425), 
      .A4(n_32_0_426), .ZN(n_32_0_427));
   AOI221_X1 i_32_0_512 (.A(n_32_0_427), .B1(\MEM[9] [5]), .B2(n_32_0_374), 
      .C1(\MEM[10] [5]), .C2(n_32_0_375), .ZN(n_32_0_428));
   AOI22_X1 i_32_0_513 (.A1(\MEM[5] [5]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [5]), .ZN(n_32_0_429));
   AOI22_X1 i_32_0_514 (.A1(\MEM[8] [5]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [5]), .ZN(n_32_0_430));
   AOI22_X1 i_32_0_515 (.A1(n_32_0_380), .A2(\MEM[6] [5]), .B1(n_32_0_381), 
      .B2(\MEM[7] [5]), .ZN(n_32_0_431));
   NAND4_X1 i_32_0_516 (.A1(n_32_0_428), .A2(n_32_0_429), .A3(n_32_0_430), 
      .A4(n_32_0_431), .ZN(data2[5]));
   AOI22_X1 i_32_0_517 (.A1(n_32_0_355), .A2(\MEM[0] [6]), .B1(n_32_0_357), 
      .B2(\MEM[2] [6]), .ZN(n_32_0_432));
   AOI22_X1 i_32_0_518 (.A1(\MEM[12] [6]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [6]), .ZN(n_32_0_433));
   AOI22_X1 i_32_0_519 (.A1(n_32_0_360), .A2(\MEM[4] [6]), .B1(n_32_0_363), 
      .B2(\MEM[13] [6]), .ZN(n_32_0_434));
   AOI22_X1 i_32_0_520 (.A1(\MEM[1] [6]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [6]), .ZN(n_32_0_435));
   NAND4_X1 i_32_0_521 (.A1(n_32_0_432), .A2(n_32_0_433), .A3(n_32_0_434), 
      .A4(n_32_0_435), .ZN(n_32_0_436));
   AOI221_X1 i_32_0_522 (.A(n_32_0_436), .B1(\MEM[9] [6]), .B2(n_32_0_374), 
      .C1(\MEM[10] [6]), .C2(n_32_0_375), .ZN(n_32_0_437));
   AOI22_X1 i_32_0_523 (.A1(\MEM[6] [6]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [6]), .ZN(n_32_0_438));
   AOI22_X1 i_32_0_524 (.A1(n_32_0_377), .A2(\MEM[8] [6]), .B1(n_32_0_378), 
      .B2(\MEM[11] [6]), .ZN(n_32_0_439));
   AOI22_X1 i_32_0_525 (.A1(\MEM[5] [6]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [6]), .ZN(n_32_0_440));
   NAND4_X1 i_32_0_526 (.A1(n_32_0_437), .A2(n_32_0_438), .A3(n_32_0_439), 
      .A4(n_32_0_440), .ZN(data2[6]));
   AOI22_X1 i_32_0_527 (.A1(n_32_0_355), .A2(\MEM[0] [7]), .B1(n_32_0_357), 
      .B2(\MEM[2] [7]), .ZN(n_32_0_441));
   AOI22_X1 i_32_0_528 (.A1(n_32_0_365), .A2(\MEM[12] [7]), .B1(n_32_0_366), 
      .B2(\MEM[14] [7]), .ZN(n_32_0_442));
   AOI22_X1 i_32_0_529 (.A1(\MEM[4] [7]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [7]), .ZN(n_32_0_443));
   AOI22_X1 i_32_0_530 (.A1(n_32_0_368), .A2(\MEM[1] [7]), .B1(n_32_0_370), 
      .B2(\MEM[15] [7]), .ZN(n_32_0_444));
   NAND4_X1 i_32_0_531 (.A1(n_32_0_441), .A2(n_32_0_442), .A3(n_32_0_443), 
      .A4(n_32_0_444), .ZN(n_32_0_445));
   AOI221_X1 i_32_0_532 (.A(n_32_0_445), .B1(\MEM[10] [7]), .B2(n_32_0_375), 
      .C1(\MEM[9] [7]), .C2(n_32_0_374), .ZN(n_32_0_446));
   AOI22_X1 i_32_0_533 (.A1(\MEM[5] [7]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [7]), .ZN(n_32_0_447));
   AOI22_X1 i_32_0_534 (.A1(n_32_0_380), .A2(\MEM[6] [7]), .B1(n_32_0_381), 
      .B2(\MEM[7] [7]), .ZN(n_32_0_448));
   AOI22_X1 i_32_0_535 (.A1(n_32_0_377), .A2(\MEM[8] [7]), .B1(n_32_0_378), 
      .B2(\MEM[11] [7]), .ZN(n_32_0_449));
   NAND4_X1 i_32_0_536 (.A1(n_32_0_446), .A2(n_32_0_447), .A3(n_32_0_448), 
      .A4(n_32_0_449), .ZN(data2[7]));
   AOI22_X1 i_32_0_537 (.A1(n_32_0_355), .A2(\MEM[0] [8]), .B1(n_32_0_357), 
      .B2(\MEM[2] [8]), .ZN(n_32_0_450));
   AOI22_X1 i_32_0_538 (.A1(\MEM[4] [8]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [8]), .ZN(n_32_0_451));
   AOI22_X1 i_32_0_539 (.A1(\MEM[12] [8]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [8]), .ZN(n_32_0_452));
   AOI22_X1 i_32_0_540 (.A1(n_32_0_368), .A2(\MEM[1] [8]), .B1(n_32_0_370), 
      .B2(\MEM[15] [8]), .ZN(n_32_0_453));
   NAND4_X1 i_32_0_541 (.A1(n_32_0_450), .A2(n_32_0_451), .A3(n_32_0_452), 
      .A4(n_32_0_453), .ZN(n_32_0_454));
   AOI221_X1 i_32_0_542 (.A(n_32_0_454), .B1(\MEM[10] [8]), .B2(n_32_0_375), 
      .C1(\MEM[9] [8]), .C2(n_32_0_374), .ZN(n_32_0_455));
   AOI22_X1 i_32_0_543 (.A1(n_32_0_383), .A2(\MEM[5] [8]), .B1(n_32_0_384), 
      .B2(\MEM[3] [8]), .ZN(n_32_0_456));
   AOI22_X1 i_32_0_544 (.A1(n_32_0_377), .A2(\MEM[8] [8]), .B1(n_32_0_378), 
      .B2(\MEM[11] [8]), .ZN(n_32_0_457));
   AOI22_X1 i_32_0_545 (.A1(\MEM[6] [8]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [8]), .ZN(n_32_0_458));
   NAND4_X1 i_32_0_546 (.A1(n_32_0_455), .A2(n_32_0_456), .A3(n_32_0_457), 
      .A4(n_32_0_458), .ZN(data2[8]));
   AOI22_X1 i_32_0_547 (.A1(n_32_0_355), .A2(\MEM[0] [9]), .B1(n_32_0_357), 
      .B2(\MEM[2] [9]), .ZN(n_32_0_459));
   AOI22_X1 i_32_0_548 (.A1(n_32_0_365), .A2(\MEM[12] [9]), .B1(n_32_0_366), 
      .B2(\MEM[14] [9]), .ZN(n_32_0_460));
   AOI22_X1 i_32_0_549 (.A1(\MEM[4] [9]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [9]), .ZN(n_32_0_461));
   AOI22_X1 i_32_0_550 (.A1(n_32_0_368), .A2(\MEM[1] [9]), .B1(n_32_0_370), 
      .B2(\MEM[15] [9]), .ZN(n_32_0_462));
   NAND4_X1 i_32_0_551 (.A1(n_32_0_459), .A2(n_32_0_460), .A3(n_32_0_461), 
      .A4(n_32_0_462), .ZN(n_32_0_463));
   AOI221_X1 i_32_0_552 (.A(n_32_0_463), .B1(\MEM[9] [9]), .B2(n_32_0_374), 
      .C1(\MEM[10] [9]), .C2(n_32_0_375), .ZN(n_32_0_464));
   AOI22_X1 i_32_0_553 (.A1(n_32_0_383), .A2(\MEM[5] [9]), .B1(n_32_0_384), 
      .B2(\MEM[3] [9]), .ZN(n_32_0_465));
   AOI22_X1 i_32_0_554 (.A1(n_32_0_377), .A2(\MEM[8] [9]), .B1(n_32_0_378), 
      .B2(\MEM[11] [9]), .ZN(n_32_0_466));
   AOI22_X1 i_32_0_555 (.A1(\MEM[6] [9]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [9]), .ZN(n_32_0_467));
   NAND4_X1 i_32_0_556 (.A1(n_32_0_464), .A2(n_32_0_465), .A3(n_32_0_466), 
      .A4(n_32_0_467), .ZN(data2[9]));
   AOI22_X1 i_32_0_557 (.A1(n_32_0_355), .A2(\MEM[0] [10]), .B1(n_32_0_357), 
      .B2(\MEM[2] [10]), .ZN(n_32_0_468));
   AOI22_X1 i_32_0_558 (.A1(n_32_0_365), .A2(\MEM[12] [10]), .B1(n_32_0_366), 
      .B2(\MEM[14] [10]), .ZN(n_32_0_469));
   AOI22_X1 i_32_0_559 (.A1(\MEM[4] [10]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [10]), .ZN(n_32_0_470));
   AOI22_X1 i_32_0_560 (.A1(n_32_0_368), .A2(\MEM[1] [10]), .B1(n_32_0_370), 
      .B2(\MEM[15] [10]), .ZN(n_32_0_471));
   NAND4_X1 i_32_0_561 (.A1(n_32_0_468), .A2(n_32_0_469), .A3(n_32_0_470), 
      .A4(n_32_0_471), .ZN(n_32_0_472));
   AOI221_X1 i_32_0_562 (.A(n_32_0_472), .B1(\MEM[9] [10]), .B2(n_32_0_374), 
      .C1(\MEM[10] [10]), .C2(n_32_0_375), .ZN(n_32_0_473));
   AOI22_X1 i_32_0_563 (.A1(n_32_0_383), .A2(\MEM[5] [10]), .B1(n_32_0_384), 
      .B2(\MEM[3] [10]), .ZN(n_32_0_474));
   AOI22_X1 i_32_0_564 (.A1(n_32_0_377), .A2(\MEM[8] [10]), .B1(n_32_0_378), 
      .B2(\MEM[11] [10]), .ZN(n_32_0_475));
   AOI22_X1 i_32_0_565 (.A1(\MEM[6] [10]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [10]), .ZN(n_32_0_476));
   NAND4_X1 i_32_0_566 (.A1(n_32_0_473), .A2(n_32_0_474), .A3(n_32_0_475), 
      .A4(n_32_0_476), .ZN(data2[10]));
   AOI22_X1 i_32_0_567 (.A1(\MEM[0] [11]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [11]), .ZN(n_32_0_477));
   AOI22_X1 i_32_0_568 (.A1(\MEM[4] [11]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [11]), .ZN(n_32_0_478));
   AOI22_X1 i_32_0_569 (.A1(\MEM[12] [11]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [11]), .ZN(n_32_0_479));
   AOI22_X1 i_32_0_570 (.A1(n_32_0_368), .A2(\MEM[1] [11]), .B1(n_32_0_370), 
      .B2(\MEM[15] [11]), .ZN(n_32_0_480));
   NAND4_X1 i_32_0_571 (.A1(n_32_0_477), .A2(n_32_0_478), .A3(n_32_0_479), 
      .A4(n_32_0_480), .ZN(n_32_0_481));
   AOI221_X1 i_32_0_572 (.A(n_32_0_481), .B1(\MEM[10] [11]), .B2(n_32_0_375), 
      .C1(\MEM[9] [11]), .C2(n_32_0_374), .ZN(n_32_0_482));
   AOI22_X1 i_32_0_573 (.A1(\MEM[5] [11]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [11]), .ZN(n_32_0_483));
   AOI22_X1 i_32_0_574 (.A1(\MEM[8] [11]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [11]), .ZN(n_32_0_484));
   AOI22_X1 i_32_0_575 (.A1(\MEM[6] [11]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [11]), .ZN(n_32_0_485));
   NAND4_X1 i_32_0_576 (.A1(n_32_0_482), .A2(n_32_0_483), .A3(n_32_0_484), 
      .A4(n_32_0_485), .ZN(data2[11]));
   AOI22_X1 i_32_0_577 (.A1(n_32_0_355), .A2(\MEM[0] [12]), .B1(n_32_0_357), 
      .B2(\MEM[2] [12]), .ZN(n_32_0_486));
   AOI22_X1 i_32_0_578 (.A1(\MEM[4] [12]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [12]), .ZN(n_32_0_487));
   AOI22_X1 i_32_0_579 (.A1(\MEM[12] [12]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [12]), .ZN(n_32_0_488));
   AOI22_X1 i_32_0_580 (.A1(\MEM[1] [12]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [12]), .ZN(n_32_0_489));
   NAND4_X1 i_32_0_581 (.A1(n_32_0_486), .A2(n_32_0_487), .A3(n_32_0_488), 
      .A4(n_32_0_489), .ZN(n_32_0_490));
   AOI221_X1 i_32_0_582 (.A(n_32_0_490), .B1(\MEM[9] [12]), .B2(n_32_0_374), 
      .C1(\MEM[10] [12]), .C2(n_32_0_375), .ZN(n_32_0_491));
   AOI22_X1 i_32_0_583 (.A1(\MEM[8] [12]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [12]), .ZN(n_32_0_492));
   AOI22_X1 i_32_0_584 (.A1(\MEM[5] [12]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [12]), .ZN(n_32_0_493));
   AOI22_X1 i_32_0_585 (.A1(\MEM[6] [12]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [12]), .ZN(n_32_0_494));
   NAND4_X1 i_32_0_586 (.A1(n_32_0_491), .A2(n_32_0_492), .A3(n_32_0_493), 
      .A4(n_32_0_494), .ZN(data2[12]));
   AOI22_X1 i_32_0_587 (.A1(n_32_0_355), .A2(\MEM[0] [13]), .B1(n_32_0_357), 
      .B2(\MEM[2] [13]), .ZN(n_32_0_495));
   AOI22_X1 i_32_0_588 (.A1(n_32_0_365), .A2(\MEM[12] [13]), .B1(n_32_0_366), 
      .B2(\MEM[14] [13]), .ZN(n_32_0_496));
   AOI22_X1 i_32_0_589 (.A1(\MEM[4] [13]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [13]), .ZN(n_32_0_497));
   AOI22_X1 i_32_0_590 (.A1(n_32_0_368), .A2(\MEM[1] [13]), .B1(n_32_0_370), 
      .B2(\MEM[15] [13]), .ZN(n_32_0_498));
   NAND4_X1 i_32_0_591 (.A1(n_32_0_495), .A2(n_32_0_496), .A3(n_32_0_497), 
      .A4(n_32_0_498), .ZN(n_32_0_499));
   AOI221_X1 i_32_0_592 (.A(n_32_0_499), .B1(\MEM[9] [13]), .B2(n_32_0_374), 
      .C1(\MEM[10] [13]), .C2(n_32_0_375), .ZN(n_32_0_500));
   AOI22_X1 i_32_0_593 (.A1(n_32_0_383), .A2(\MEM[5] [13]), .B1(n_32_0_384), 
      .B2(\MEM[3] [13]), .ZN(n_32_0_501));
   AOI22_X1 i_32_0_594 (.A1(n_32_0_377), .A2(\MEM[8] [13]), .B1(n_32_0_378), 
      .B2(\MEM[11] [13]), .ZN(n_32_0_502));
   AOI22_X1 i_32_0_595 (.A1(\MEM[6] [13]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [13]), .ZN(n_32_0_503));
   NAND4_X1 i_32_0_596 (.A1(n_32_0_500), .A2(n_32_0_501), .A3(n_32_0_502), 
      .A4(n_32_0_503), .ZN(data2[13]));
   AOI22_X1 i_32_0_597 (.A1(n_32_0_355), .A2(\MEM[0] [14]), .B1(n_32_0_357), 
      .B2(\MEM[2] [14]), .ZN(n_32_0_504));
   AOI22_X1 i_32_0_598 (.A1(n_32_0_360), .A2(\MEM[4] [14]), .B1(n_32_0_363), 
      .B2(\MEM[13] [14]), .ZN(n_32_0_505));
   AOI22_X1 i_32_0_599 (.A1(\MEM[12] [14]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [14]), .ZN(n_32_0_506));
   AOI22_X1 i_32_0_600 (.A1(n_32_0_368), .A2(\MEM[1] [14]), .B1(n_32_0_370), 
      .B2(\MEM[15] [14]), .ZN(n_32_0_507));
   NAND4_X1 i_32_0_601 (.A1(n_32_0_504), .A2(n_32_0_505), .A3(n_32_0_506), 
      .A4(n_32_0_507), .ZN(n_32_0_508));
   AOI221_X1 i_32_0_602 (.A(n_32_0_508), .B1(\MEM[10] [14]), .B2(n_32_0_375), 
      .C1(\MEM[9] [14]), .C2(n_32_0_374), .ZN(n_32_0_509));
   AOI22_X1 i_32_0_603 (.A1(n_32_0_377), .A2(\MEM[8] [14]), .B1(n_32_0_378), 
      .B2(\MEM[11] [14]), .ZN(n_32_0_510));
   AOI22_X1 i_32_0_604 (.A1(n_32_0_383), .A2(\MEM[5] [14]), .B1(n_32_0_384), 
      .B2(\MEM[3] [14]), .ZN(n_32_0_511));
   AOI22_X1 i_32_0_605 (.A1(n_32_0_380), .A2(\MEM[6] [14]), .B1(n_32_0_381), 
      .B2(\MEM[7] [14]), .ZN(n_32_0_512));
   NAND4_X1 i_32_0_606 (.A1(n_32_0_509), .A2(n_32_0_510), .A3(n_32_0_511), 
      .A4(n_32_0_512), .ZN(data2[14]));
   AOI22_X1 i_32_0_607 (.A1(n_32_0_355), .A2(\MEM[0] [15]), .B1(n_32_0_357), 
      .B2(\MEM[2] [15]), .ZN(n_32_0_513));
   AOI22_X1 i_32_0_608 (.A1(n_32_0_365), .A2(\MEM[12] [15]), .B1(n_32_0_366), 
      .B2(\MEM[14] [15]), .ZN(n_32_0_514));
   AOI22_X1 i_32_0_609 (.A1(\MEM[4] [15]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [15]), .ZN(n_32_0_515));
   AOI22_X1 i_32_0_610 (.A1(n_32_0_368), .A2(\MEM[1] [15]), .B1(n_32_0_370), 
      .B2(\MEM[15] [15]), .ZN(n_32_0_516));
   NAND4_X1 i_32_0_611 (.A1(n_32_0_513), .A2(n_32_0_514), .A3(n_32_0_515), 
      .A4(n_32_0_516), .ZN(n_32_0_517));
   AOI221_X1 i_32_0_612 (.A(n_32_0_517), .B1(\MEM[9] [15]), .B2(n_32_0_374), 
      .C1(\MEM[10] [15]), .C2(n_32_0_375), .ZN(n_32_0_518));
   AOI22_X1 i_32_0_613 (.A1(n_32_0_383), .A2(\MEM[5] [15]), .B1(n_32_0_384), 
      .B2(\MEM[3] [15]), .ZN(n_32_0_519));
   AOI22_X1 i_32_0_614 (.A1(n_32_0_377), .A2(\MEM[8] [15]), .B1(n_32_0_378), 
      .B2(\MEM[11] [15]), .ZN(n_32_0_520));
   AOI22_X1 i_32_0_615 (.A1(\MEM[6] [15]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [15]), .ZN(n_32_0_521));
   NAND4_X1 i_32_0_616 (.A1(n_32_0_518), .A2(n_32_0_519), .A3(n_32_0_520), 
      .A4(n_32_0_521), .ZN(data2[15]));
   AOI22_X1 i_32_0_617 (.A1(n_32_0_355), .A2(\MEM[0] [16]), .B1(n_32_0_357), 
      .B2(\MEM[2] [16]), .ZN(n_32_0_522));
   AOI22_X1 i_32_0_618 (.A1(\MEM[4] [16]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [16]), .ZN(n_32_0_523));
   AOI22_X1 i_32_0_619 (.A1(n_32_0_365), .A2(\MEM[12] [16]), .B1(n_32_0_366), 
      .B2(\MEM[14] [16]), .ZN(n_32_0_524));
   AOI22_X1 i_32_0_620 (.A1(n_32_0_368), .A2(\MEM[1] [16]), .B1(n_32_0_370), 
      .B2(\MEM[15] [16]), .ZN(n_32_0_525));
   NAND4_X1 i_32_0_621 (.A1(n_32_0_522), .A2(n_32_0_523), .A3(n_32_0_524), 
      .A4(n_32_0_525), .ZN(n_32_0_526));
   AOI221_X1 i_32_0_622 (.A(n_32_0_526), .B1(\MEM[9] [16]), .B2(n_32_0_374), 
      .C1(\MEM[10] [16]), .C2(n_32_0_375), .ZN(n_32_0_527));
   AOI22_X1 i_32_0_623 (.A1(\MEM[8] [16]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [16]), .ZN(n_32_0_528));
   AOI22_X1 i_32_0_624 (.A1(\MEM[5] [16]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [16]), .ZN(n_32_0_529));
   AOI22_X1 i_32_0_625 (.A1(\MEM[6] [16]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [16]), .ZN(n_32_0_530));
   NAND4_X1 i_32_0_626 (.A1(n_32_0_527), .A2(n_32_0_528), .A3(n_32_0_529), 
      .A4(n_32_0_530), .ZN(data2[16]));
   AOI22_X1 i_32_0_627 (.A1(n_32_0_355), .A2(\MEM[0] [17]), .B1(n_32_0_357), 
      .B2(\MEM[2] [17]), .ZN(n_32_0_531));
   AOI22_X1 i_32_0_628 (.A1(\MEM[12] [17]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [17]), .ZN(n_32_0_532));
   AOI22_X1 i_32_0_629 (.A1(\MEM[4] [17]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [17]), .ZN(n_32_0_533));
   AOI22_X1 i_32_0_630 (.A1(n_32_0_368), .A2(\MEM[1] [17]), .B1(n_32_0_370), 
      .B2(\MEM[15] [17]), .ZN(n_32_0_534));
   NAND4_X1 i_32_0_631 (.A1(n_32_0_531), .A2(n_32_0_532), .A3(n_32_0_533), 
      .A4(n_32_0_534), .ZN(n_32_0_535));
   AOI221_X1 i_32_0_632 (.A(n_32_0_535), .B1(\MEM[9] [17]), .B2(n_32_0_374), 
      .C1(\MEM[10] [17]), .C2(n_32_0_375), .ZN(n_32_0_536));
   AOI22_X1 i_32_0_633 (.A1(n_32_0_383), .A2(\MEM[5] [17]), .B1(n_32_0_384), 
      .B2(\MEM[3] [17]), .ZN(n_32_0_537));
   AOI22_X1 i_32_0_634 (.A1(n_32_0_377), .A2(\MEM[8] [17]), .B1(n_32_0_378), 
      .B2(\MEM[11] [17]), .ZN(n_32_0_538));
   AOI22_X1 i_32_0_635 (.A1(\MEM[6] [17]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [17]), .ZN(n_32_0_539));
   NAND4_X1 i_32_0_636 (.A1(n_32_0_536), .A2(n_32_0_537), .A3(n_32_0_538), 
      .A4(n_32_0_539), .ZN(data2[17]));
   AOI22_X1 i_32_0_637 (.A1(\MEM[0] [18]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [18]), .ZN(n_32_0_540));
   AOI22_X1 i_32_0_638 (.A1(\MEM[12] [18]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [18]), .ZN(n_32_0_541));
   AOI22_X1 i_32_0_639 (.A1(\MEM[4] [18]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [18]), .ZN(n_32_0_542));
   AOI22_X1 i_32_0_640 (.A1(n_32_0_368), .A2(\MEM[1] [18]), .B1(n_32_0_370), 
      .B2(\MEM[15] [18]), .ZN(n_32_0_543));
   NAND4_X1 i_32_0_641 (.A1(n_32_0_540), .A2(n_32_0_541), .A3(n_32_0_542), 
      .A4(n_32_0_543), .ZN(n_32_0_544));
   AOI221_X1 i_32_0_642 (.A(n_32_0_544), .B1(\MEM[9] [18]), .B2(n_32_0_374), 
      .C1(\MEM[10] [18]), .C2(n_32_0_375), .ZN(n_32_0_545));
   AOI22_X1 i_32_0_643 (.A1(n_32_0_380), .A2(\MEM[6] [18]), .B1(n_32_0_381), 
      .B2(\MEM[7] [18]), .ZN(n_32_0_546));
   AOI22_X1 i_32_0_644 (.A1(\MEM[8] [18]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [18]), .ZN(n_32_0_547));
   AOI22_X1 i_32_0_645 (.A1(\MEM[5] [18]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [18]), .ZN(n_32_0_548));
   NAND4_X1 i_32_0_646 (.A1(n_32_0_545), .A2(n_32_0_546), .A3(n_32_0_547), 
      .A4(n_32_0_548), .ZN(data2[18]));
   AOI22_X1 i_32_0_647 (.A1(\MEM[6] [19]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [19]), .ZN(n_32_0_549));
   AOI22_X1 i_32_0_648 (.A1(n_32_0_377), .A2(\MEM[8] [19]), .B1(n_32_0_378), 
      .B2(\MEM[11] [19]), .ZN(n_32_0_550));
   NAND2_X1 i_32_0_649 (.A1(n_32_0_549), .A2(n_32_0_550), .ZN(n_32_0_551));
   AOI221_X1 i_32_0_650 (.A(n_32_0_551), .B1(\MEM[3] [19]), .B2(n_32_0_384), 
      .C1(\MEM[5] [19]), .C2(n_32_0_383), .ZN(n_32_0_552));
   AOI22_X1 i_32_0_651 (.A1(\MEM[12] [19]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [19]), .ZN(n_32_0_553));
   AOI22_X1 i_32_0_652 (.A1(\MEM[1] [19]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [19]), .ZN(n_32_0_554));
   NAND2_X1 i_32_0_653 (.A1(n_32_0_553), .A2(n_32_0_554), .ZN(n_32_0_555));
   AOI221_X1 i_32_0_654 (.A(n_32_0_555), .B1(\MEM[13] [19]), .B2(n_32_0_363), 
      .C1(\MEM[4] [19]), .C2(n_32_0_360), .ZN(n_32_0_556));
   AOI22_X1 i_32_0_655 (.A1(\MEM[0] [19]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [19]), .ZN(n_32_0_557));
   AOI22_X1 i_32_0_656 (.A1(n_32_0_374), .A2(\MEM[9] [19]), .B1(n_32_0_375), 
      .B2(\MEM[10] [19]), .ZN(n_32_0_558));
   NAND4_X1 i_32_0_657 (.A1(n_32_0_552), .A2(n_32_0_556), .A3(n_32_0_557), 
      .A4(n_32_0_558), .ZN(data2[19]));
   AOI22_X1 i_32_0_658 (.A1(n_32_0_355), .A2(\MEM[0] [20]), .B1(n_32_0_357), 
      .B2(\MEM[2] [20]), .ZN(n_32_0_559));
   AOI22_X1 i_32_0_659 (.A1(n_32_0_360), .A2(\MEM[4] [20]), .B1(n_32_0_363), 
      .B2(\MEM[13] [20]), .ZN(n_32_0_560));
   AOI22_X1 i_32_0_660 (.A1(\MEM[12] [20]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [20]), .ZN(n_32_0_561));
   AOI22_X1 i_32_0_661 (.A1(n_32_0_368), .A2(\MEM[1] [20]), .B1(n_32_0_370), 
      .B2(\MEM[15] [20]), .ZN(n_32_0_562));
   NAND4_X1 i_32_0_662 (.A1(n_32_0_559), .A2(n_32_0_560), .A3(n_32_0_561), 
      .A4(n_32_0_562), .ZN(n_32_0_563));
   AOI221_X1 i_32_0_663 (.A(n_32_0_563), .B1(\MEM[10] [20]), .B2(n_32_0_375), 
      .C1(\MEM[9] [20]), .C2(n_32_0_374), .ZN(n_32_0_564));
   AOI22_X1 i_32_0_664 (.A1(\MEM[5] [20]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [20]), .ZN(n_32_0_565));
   AOI22_X1 i_32_0_665 (.A1(n_32_0_380), .A2(\MEM[6] [20]), .B1(n_32_0_381), 
      .B2(\MEM[7] [20]), .ZN(n_32_0_566));
   AOI22_X1 i_32_0_666 (.A1(n_32_0_377), .A2(\MEM[8] [20]), .B1(n_32_0_378), 
      .B2(\MEM[11] [20]), .ZN(n_32_0_567));
   NAND4_X1 i_32_0_667 (.A1(n_32_0_564), .A2(n_32_0_565), .A3(n_32_0_566), 
      .A4(n_32_0_567), .ZN(data2[20]));
   AOI22_X1 i_32_0_668 (.A1(\MEM[0] [21]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [21]), .ZN(n_32_0_568));
   AOI22_X1 i_32_0_669 (.A1(n_32_0_365), .A2(\MEM[12] [21]), .B1(n_32_0_366), 
      .B2(\MEM[14] [21]), .ZN(n_32_0_569));
   NAND2_X1 i_32_0_670 (.A1(n_32_0_568), .A2(n_32_0_569), .ZN(n_32_0_570));
   AOI221_X1 i_32_0_671 (.A(n_32_0_570), .B1(\MEM[13] [21]), .B2(n_32_0_363), 
      .C1(\MEM[4] [21]), .C2(n_32_0_360), .ZN(n_32_0_571));
   AOI22_X1 i_32_0_672 (.A1(\MEM[5] [21]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [21]), .ZN(n_32_0_572));
   AOI22_X1 i_32_0_673 (.A1(n_32_0_380), .A2(\MEM[6] [21]), .B1(n_32_0_381), 
      .B2(\MEM[7] [21]), .ZN(n_32_0_573));
   NAND2_X1 i_32_0_674 (.A1(n_32_0_572), .A2(n_32_0_573), .ZN(n_32_0_574));
   AOI221_X1 i_32_0_675 (.A(n_32_0_574), .B1(\MEM[11] [21]), .B2(n_32_0_378), 
      .C1(\MEM[8] [21]), .C2(n_32_0_377), .ZN(n_32_0_575));
   AOI22_X1 i_32_0_676 (.A1(\MEM[1] [21]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [21]), .ZN(n_32_0_576));
   AOI22_X1 i_32_0_677 (.A1(n_32_0_375), .A2(\MEM[10] [21]), .B1(n_32_0_374), 
      .B2(\MEM[9] [21]), .ZN(n_32_0_577));
   NAND4_X1 i_32_0_678 (.A1(n_32_0_571), .A2(n_32_0_575), .A3(n_32_0_576), 
      .A4(n_32_0_577), .ZN(data2[21]));
   AOI22_X1 i_32_0_679 (.A1(n_32_0_355), .A2(\MEM[0] [22]), .B1(n_32_0_357), 
      .B2(\MEM[2] [22]), .ZN(n_32_0_578));
   AOI22_X1 i_32_0_680 (.A1(n_32_0_360), .A2(\MEM[4] [22]), .B1(n_32_0_363), 
      .B2(\MEM[13] [22]), .ZN(n_32_0_579));
   AOI22_X1 i_32_0_681 (.A1(n_32_0_365), .A2(\MEM[12] [22]), .B1(n_32_0_366), 
      .B2(\MEM[14] [22]), .ZN(n_32_0_580));
   AOI22_X1 i_32_0_682 (.A1(n_32_0_368), .A2(\MEM[1] [22]), .B1(n_32_0_370), 
      .B2(\MEM[15] [22]), .ZN(n_32_0_581));
   NAND4_X1 i_32_0_683 (.A1(n_32_0_578), .A2(n_32_0_579), .A3(n_32_0_580), 
      .A4(n_32_0_581), .ZN(n_32_0_582));
   AOI221_X1 i_32_0_684 (.A(n_32_0_582), .B1(\MEM[10] [22]), .B2(n_32_0_375), 
      .C1(\MEM[9] [22]), .C2(n_32_0_374), .ZN(n_32_0_583));
   AOI22_X1 i_32_0_685 (.A1(\MEM[5] [22]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [22]), .ZN(n_32_0_584));
   AOI22_X1 i_32_0_686 (.A1(n_32_0_380), .A2(\MEM[6] [22]), .B1(n_32_0_381), 
      .B2(\MEM[7] [22]), .ZN(n_32_0_585));
   AOI22_X1 i_32_0_687 (.A1(\MEM[8] [22]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [22]), .ZN(n_32_0_586));
   NAND4_X1 i_32_0_688 (.A1(n_32_0_583), .A2(n_32_0_584), .A3(n_32_0_585), 
      .A4(n_32_0_586), .ZN(data2[22]));
   AOI22_X1 i_32_0_689 (.A1(n_32_0_355), .A2(\MEM[0] [23]), .B1(n_32_0_357), 
      .B2(\MEM[2] [23]), .ZN(n_32_0_587));
   AOI22_X1 i_32_0_690 (.A1(\MEM[12] [23]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [23]), .ZN(n_32_0_588));
   AOI22_X1 i_32_0_691 (.A1(n_32_0_360), .A2(\MEM[4] [23]), .B1(n_32_0_363), 
      .B2(\MEM[13] [23]), .ZN(n_32_0_589));
   AOI22_X1 i_32_0_692 (.A1(n_32_0_368), .A2(\MEM[1] [23]), .B1(n_32_0_370), 
      .B2(\MEM[15] [23]), .ZN(n_32_0_590));
   NAND4_X1 i_32_0_693 (.A1(n_32_0_587), .A2(n_32_0_588), .A3(n_32_0_589), 
      .A4(n_32_0_590), .ZN(n_32_0_591));
   AOI221_X1 i_32_0_694 (.A(n_32_0_591), .B1(\MEM[10] [23]), .B2(n_32_0_375), 
      .C1(\MEM[9] [23]), .C2(n_32_0_374), .ZN(n_32_0_592));
   AOI22_X1 i_32_0_695 (.A1(\MEM[5] [23]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [23]), .ZN(n_32_0_593));
   AOI22_X1 i_32_0_696 (.A1(n_32_0_380), .A2(\MEM[6] [23]), .B1(n_32_0_381), 
      .B2(\MEM[7] [23]), .ZN(n_32_0_594));
   AOI22_X1 i_32_0_697 (.A1(n_32_0_377), .A2(\MEM[8] [23]), .B1(n_32_0_378), 
      .B2(\MEM[11] [23]), .ZN(n_32_0_595));
   NAND4_X1 i_32_0_698 (.A1(n_32_0_592), .A2(n_32_0_593), .A3(n_32_0_594), 
      .A4(n_32_0_595), .ZN(data2[23]));
   AOI22_X1 i_32_0_699 (.A1(n_32_0_355), .A2(\MEM[0] [24]), .B1(n_32_0_357), 
      .B2(\MEM[2] [24]), .ZN(n_32_0_596));
   AOI22_X1 i_32_0_700 (.A1(n_32_0_365), .A2(\MEM[12] [24]), .B1(n_32_0_366), 
      .B2(\MEM[14] [24]), .ZN(n_32_0_597));
   AOI22_X1 i_32_0_701 (.A1(n_32_0_360), .A2(\MEM[4] [24]), .B1(n_32_0_363), 
      .B2(\MEM[13] [24]), .ZN(n_32_0_598));
   AOI22_X1 i_32_0_702 (.A1(n_32_0_368), .A2(\MEM[1] [24]), .B1(n_32_0_370), 
      .B2(\MEM[15] [24]), .ZN(n_32_0_599));
   NAND4_X1 i_32_0_703 (.A1(n_32_0_596), .A2(n_32_0_597), .A3(n_32_0_598), 
      .A4(n_32_0_599), .ZN(n_32_0_600));
   AOI221_X1 i_32_0_704 (.A(n_32_0_600), .B1(\MEM[10] [24]), .B2(n_32_0_375), 
      .C1(\MEM[9] [24]), .C2(n_32_0_374), .ZN(n_32_0_601));
   AOI22_X1 i_32_0_705 (.A1(n_32_0_380), .A2(\MEM[6] [24]), .B1(n_32_0_381), 
      .B2(\MEM[7] [24]), .ZN(n_32_0_602));
   AOI22_X1 i_32_0_706 (.A1(\MEM[8] [24]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [24]), .ZN(n_32_0_603));
   AOI22_X1 i_32_0_707 (.A1(\MEM[5] [24]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [24]), .ZN(n_32_0_604));
   NAND4_X1 i_32_0_708 (.A1(n_32_0_601), .A2(n_32_0_602), .A3(n_32_0_603), 
      .A4(n_32_0_604), .ZN(data2[24]));
   AOI22_X1 i_32_0_709 (.A1(n_32_0_355), .A2(\MEM[0] [25]), .B1(n_32_0_357), 
      .B2(\MEM[2] [25]), .ZN(n_32_0_605));
   AOI22_X1 i_32_0_710 (.A1(\MEM[12] [25]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [25]), .ZN(n_32_0_606));
   AOI22_X1 i_32_0_711 (.A1(\MEM[4] [25]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [25]), .ZN(n_32_0_607));
   AOI22_X1 i_32_0_712 (.A1(n_32_0_368), .A2(\MEM[1] [25]), .B1(n_32_0_370), 
      .B2(\MEM[15] [25]), .ZN(n_32_0_608));
   NAND4_X1 i_32_0_713 (.A1(n_32_0_605), .A2(n_32_0_606), .A3(n_32_0_607), 
      .A4(n_32_0_608), .ZN(n_32_0_609));
   AOI221_X1 i_32_0_714 (.A(n_32_0_609), .B1(\MEM[9] [25]), .B2(n_32_0_374), 
      .C1(\MEM[10] [25]), .C2(n_32_0_375), .ZN(n_32_0_610));
   AOI22_X1 i_32_0_715 (.A1(\MEM[5] [25]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [25]), .ZN(n_32_0_611));
   AOI22_X1 i_32_0_716 (.A1(n_32_0_377), .A2(\MEM[8] [25]), .B1(n_32_0_378), 
      .B2(\MEM[11] [25]), .ZN(n_32_0_612));
   AOI22_X1 i_32_0_717 (.A1(n_32_0_380), .A2(\MEM[6] [25]), .B1(n_32_0_381), 
      .B2(\MEM[7] [25]), .ZN(n_32_0_613));
   NAND4_X1 i_32_0_718 (.A1(n_32_0_610), .A2(n_32_0_611), .A3(n_32_0_612), 
      .A4(n_32_0_613), .ZN(data2[25]));
   AOI22_X1 i_32_0_719 (.A1(\MEM[0] [26]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [26]), .ZN(n_32_0_614));
   AOI22_X1 i_32_0_720 (.A1(n_32_0_360), .A2(\MEM[4] [26]), .B1(n_32_0_363), 
      .B2(\MEM[13] [26]), .ZN(n_32_0_615));
   NAND2_X1 i_32_0_721 (.A1(n_32_0_614), .A2(n_32_0_615), .ZN(n_32_0_616));
   AOI221_X1 i_32_0_722 (.A(n_32_0_616), .B1(\MEM[14] [26]), .B2(n_32_0_366), 
      .C1(\MEM[12] [26]), .C2(n_32_0_365), .ZN(n_32_0_617));
   AOI22_X1 i_32_0_723 (.A1(\MEM[8] [26]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [26]), .ZN(n_32_0_618));
   AOI22_X1 i_32_0_724 (.A1(n_32_0_380), .A2(\MEM[6] [26]), .B1(n_32_0_381), 
      .B2(\MEM[7] [26]), .ZN(n_32_0_619));
   NAND2_X1 i_32_0_725 (.A1(n_32_0_618), .A2(n_32_0_619), .ZN(n_32_0_620));
   AOI221_X1 i_32_0_726 (.A(n_32_0_620), .B1(\MEM[3] [26]), .B2(n_32_0_384), 
      .C1(\MEM[5] [26]), .C2(n_32_0_383), .ZN(n_32_0_621));
   AOI22_X1 i_32_0_727 (.A1(\MEM[1] [26]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [26]), .ZN(n_32_0_622));
   AOI22_X1 i_32_0_728 (.A1(n_32_0_375), .A2(\MEM[10] [26]), .B1(n_32_0_374), 
      .B2(\MEM[9] [26]), .ZN(n_32_0_623));
   NAND4_X1 i_32_0_729 (.A1(n_32_0_617), .A2(n_32_0_621), .A3(n_32_0_622), 
      .A4(n_32_0_623), .ZN(data2[26]));
   AOI22_X1 i_32_0_730 (.A1(\MEM[0] [27]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [27]), .ZN(n_32_0_624));
   AOI22_X1 i_32_0_731 (.A1(n_32_0_360), .A2(\MEM[4] [27]), .B1(n_32_0_363), 
      .B2(\MEM[13] [27]), .ZN(n_32_0_625));
   AOI22_X1 i_32_0_732 (.A1(\MEM[1] [27]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [27]), .ZN(n_32_0_626));
   NAND3_X1 i_32_0_733 (.A1(n_32_0_624), .A2(n_32_0_625), .A3(n_32_0_626), 
      .ZN(n_32_0_627));
   AOI221_X1 i_32_0_734 (.A(n_32_0_627), .B1(\MEM[12] [27]), .B2(n_32_0_365), 
      .C1(\MEM[14] [27]), .C2(n_32_0_366), .ZN(n_32_0_628));
   AOI222_X1 i_32_0_735 (.A1(n_32_0_375), .A2(\MEM[10] [27]), .B1(n_32_0_374), 
      .B2(\MEM[9] [27]), .C1(n_32_0_384), .C2(\MEM[3] [27]), .ZN(n_32_0_629));
   AOI22_X1 i_32_0_736 (.A1(\MEM[8] [27]), .A2(n_32_0_377), .B1(n_32_0_383), 
      .B2(\MEM[5] [27]), .ZN(n_32_0_630));
   AOI222_X1 i_32_0_737 (.A1(n_32_0_380), .A2(\MEM[6] [27]), .B1(n_32_0_381), 
      .B2(\MEM[7] [27]), .C1(n_32_0_378), .C2(\MEM[11] [27]), .ZN(n_32_0_631));
   NAND4_X1 i_32_0_738 (.A1(n_32_0_628), .A2(n_32_0_629), .A3(n_32_0_630), 
      .A4(n_32_0_631), .ZN(data2[27]));
   AOI22_X1 i_32_0_739 (.A1(n_32_0_355), .A2(\MEM[0] [28]), .B1(n_32_0_357), 
      .B2(\MEM[2] [28]), .ZN(n_32_0_632));
   AOI22_X1 i_32_0_740 (.A1(\MEM[12] [28]), .A2(n_32_0_365), .B1(n_32_0_366), 
      .B2(\MEM[14] [28]), .ZN(n_32_0_633));
   AOI22_X1 i_32_0_741 (.A1(\MEM[4] [28]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [28]), .ZN(n_32_0_634));
   AOI22_X1 i_32_0_742 (.A1(\MEM[1] [28]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [28]), .ZN(n_32_0_635));
   NAND4_X1 i_32_0_743 (.A1(n_32_0_632), .A2(n_32_0_633), .A3(n_32_0_634), 
      .A4(n_32_0_635), .ZN(n_32_0_636));
   AOI221_X1 i_32_0_744 (.A(n_32_0_636), .B1(\MEM[9] [28]), .B2(n_32_0_374), 
      .C1(\MEM[10] [28]), .C2(n_32_0_375), .ZN(n_32_0_637));
   AOI22_X1 i_32_0_745 (.A1(\MEM[6] [28]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [28]), .ZN(n_32_0_638));
   AOI22_X1 i_32_0_746 (.A1(\MEM[8] [28]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [28]), .ZN(n_32_0_639));
   AOI22_X1 i_32_0_747 (.A1(\MEM[5] [28]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [28]), .ZN(n_32_0_640));
   NAND4_X1 i_32_0_748 (.A1(n_32_0_637), .A2(n_32_0_638), .A3(n_32_0_639), 
      .A4(n_32_0_640), .ZN(data2[28]));
   AOI22_X1 i_32_0_749 (.A1(n_32_0_355), .A2(\MEM[0] [29]), .B1(n_32_0_357), 
      .B2(\MEM[2] [29]), .ZN(n_32_0_641));
   AOI22_X1 i_32_0_750 (.A1(n_32_0_365), .A2(\MEM[12] [29]), .B1(n_32_0_366), 
      .B2(\MEM[14] [29]), .ZN(n_32_0_642));
   AOI22_X1 i_32_0_751 (.A1(\MEM[4] [29]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [29]), .ZN(n_32_0_643));
   AOI22_X1 i_32_0_752 (.A1(n_32_0_368), .A2(\MEM[1] [29]), .B1(n_32_0_370), 
      .B2(\MEM[15] [29]), .ZN(n_32_0_644));
   NAND4_X1 i_32_0_753 (.A1(n_32_0_641), .A2(n_32_0_642), .A3(n_32_0_643), 
      .A4(n_32_0_644), .ZN(n_32_0_645));
   AOI221_X1 i_32_0_754 (.A(n_32_0_645), .B1(\MEM[9] [29]), .B2(n_32_0_374), 
      .C1(\MEM[10] [29]), .C2(n_32_0_375), .ZN(n_32_0_646));
   AOI22_X1 i_32_0_755 (.A1(n_32_0_383), .A2(\MEM[5] [29]), .B1(n_32_0_384), 
      .B2(\MEM[3] [29]), .ZN(n_32_0_647));
   AOI22_X1 i_32_0_756 (.A1(n_32_0_377), .A2(\MEM[8] [29]), .B1(n_32_0_378), 
      .B2(\MEM[11] [29]), .ZN(n_32_0_648));
   AOI22_X1 i_32_0_757 (.A1(\MEM[6] [29]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [29]), .ZN(n_32_0_649));
   NAND4_X1 i_32_0_758 (.A1(n_32_0_646), .A2(n_32_0_647), .A3(n_32_0_648), 
      .A4(n_32_0_649), .ZN(data2[29]));
   AOI22_X1 i_32_0_759 (.A1(\MEM[0] [30]), .A2(n_32_0_355), .B1(n_32_0_357), 
      .B2(\MEM[2] [30]), .ZN(n_32_0_650));
   AOI22_X1 i_32_0_760 (.A1(n_32_0_365), .A2(\MEM[12] [30]), .B1(n_32_0_366), 
      .B2(\MEM[14] [30]), .ZN(n_32_0_651));
   AOI22_X1 i_32_0_761 (.A1(\MEM[4] [30]), .A2(n_32_0_360), .B1(n_32_0_363), 
      .B2(\MEM[13] [30]), .ZN(n_32_0_652));
   AOI22_X1 i_32_0_762 (.A1(n_32_0_368), .A2(\MEM[1] [30]), .B1(n_32_0_370), 
      .B2(\MEM[15] [30]), .ZN(n_32_0_653));
   NAND4_X1 i_32_0_763 (.A1(n_32_0_650), .A2(n_32_0_651), .A3(n_32_0_652), 
      .A4(n_32_0_653), .ZN(n_32_0_654));
   AOI221_X1 i_32_0_764 (.A(n_32_0_654), .B1(\MEM[10] [30]), .B2(n_32_0_375), 
      .C1(\MEM[9] [30]), .C2(n_32_0_374), .ZN(n_32_0_655));
   AOI22_X1 i_32_0_765 (.A1(\MEM[8] [30]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [30]), .ZN(n_32_0_656));
   AOI22_X1 i_32_0_766 (.A1(n_32_0_380), .A2(\MEM[6] [30]), .B1(n_32_0_381), 
      .B2(\MEM[7] [30]), .ZN(n_32_0_657));
   AOI22_X1 i_32_0_767 (.A1(\MEM[5] [30]), .A2(n_32_0_383), .B1(n_32_0_384), 
      .B2(\MEM[3] [30]), .ZN(n_32_0_658));
   NAND4_X1 i_32_0_768 (.A1(n_32_0_655), .A2(n_32_0_656), .A3(n_32_0_657), 
      .A4(n_32_0_658), .ZN(data2[30]));
   AOI22_X1 i_32_0_769 (.A1(n_32_0_365), .A2(\MEM[12] [31]), .B1(n_32_0_363), 
      .B2(\MEM[13] [31]), .ZN(n_32_0_659));
   AOI22_X1 i_32_0_770 (.A1(n_32_0_360), .A2(\MEM[4] [31]), .B1(n_32_0_384), 
      .B2(\MEM[3] [31]), .ZN(n_32_0_660));
   AOI22_X1 i_32_0_771 (.A1(n_32_0_355), .A2(\MEM[0] [31]), .B1(n_32_0_366), 
      .B2(\MEM[14] [31]), .ZN(n_32_0_661));
   AOI22_X1 i_32_0_772 (.A1(\MEM[1] [31]), .A2(n_32_0_368), .B1(n_32_0_370), 
      .B2(\MEM[15] [31]), .ZN(n_32_0_662));
   NAND4_X1 i_32_0_773 (.A1(n_32_0_659), .A2(n_32_0_660), .A3(n_32_0_661), 
      .A4(n_32_0_662), .ZN(n_32_0_663));
   AOI221_X1 i_32_0_774 (.A(n_32_0_663), .B1(\MEM[10] [31]), .B2(n_32_0_375), 
      .C1(\MEM[9] [31]), .C2(n_32_0_374), .ZN(n_32_0_664));
   AOI22_X1 i_32_0_775 (.A1(n_32_0_357), .A2(\MEM[2] [31]), .B1(n_32_0_383), 
      .B2(\MEM[5] [31]), .ZN(n_32_0_665));
   AOI22_X1 i_32_0_776 (.A1(\MEM[6] [31]), .A2(n_32_0_380), .B1(n_32_0_381), 
      .B2(\MEM[7] [31]), .ZN(n_32_0_666));
   AOI22_X1 i_32_0_777 (.A1(\MEM[8] [31]), .A2(n_32_0_377), .B1(n_32_0_378), 
      .B2(\MEM[11] [31]), .ZN(n_32_0_667));
   NAND4_X1 i_32_0_778 (.A1(n_32_0_664), .A2(n_32_0_665), .A3(n_32_0_666), 
      .A4(n_32_0_667), .ZN(data2[31]));
   INV_X1 i_32_0_779 (.A(n_32_0_348), .ZN(MEM[31]));
endmodule
