module MAIN_EULAR (
);


endmodule