/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Apr 23 16:55:22 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3334430703 */

module multiplier(clk, rst, multiplicand, multiplier, start, result, 
      overflow_flag, finish);
   input clk;
   input rst;
   input [15:0]multiplicand;
   input [15:0]multiplier;
   input start;
   output [15:0]result;
   output overflow_flag;
   output finish;

   wire n_0_2;
   wire [15:0]A;
   wire n_0_0;
   wire [15:0]multiplicand_buffer;
   wire [16:0]Q;
   wire [2:0]counter;
   wire working;
   wire start_buffer;
   wire n_0_3;
   wire n_0_1;
   wire n_0_6;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_7;
   wire n_0_0_2;
   wire n_0_8;
   wire n_0_0_3;
   wire n_0_9;
   wire n_0_0_5;
   wire n_0_10;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_12;
   wire n_0_18;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_19;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_32;
   wire n_0_0_64;
   wire n_0_0_17;
   wire n_0_0_69;
   wire n_0_0_18;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_20;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_21;
   wire n_0_22;
   wire n_0_0_148;
   wire n_0_23;
   wire n_0_0_149;
   wire n_0_24;
   wire n_0_0_150;
   wire n_0_25;
   wire n_0_0_151;
   wire n_0_26;
   wire n_0_0_152;
   wire n_0_27;
   wire n_0_0_153;
   wire n_0_28;
   wire n_0_0_154;
   wire n_0_29;
   wire n_0_0_155;
   wire n_0_30;
   wire n_0_0_156;
   wire n_0_31;
   wire n_0_0_157;
   wire n_0_32;
   wire n_0_0_158;
   wire n_0_33;
   wire n_0_0_159;
   wire n_0_34;
   wire n_0_0_160;
   wire n_0_35;
   wire n_0_0_161;
   wire n_0_36;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_37;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_19;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_20;
   wire n_0_0_171;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_38;
   wire n_0_4;
   wire n_0_39;
   wire n_0_40;
   wire n_0_0_184;
   wire n_0_41;
   wire n_0_0_185;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_60;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_4;
   wire n_0_0_6;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_21;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_5;
   wire n_0_0_22;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_11;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_13;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_14;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_15;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_59;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_16;
   wire n_0_0_137;
   wire n_0_17;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_167;
   wire n_0_0_170;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_178;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_186;
   wire n_0_0_187;

   INV_X1 adder_counter_which_adder_0_adder_block_inst1_full_adder_inst1_i_3 (
      .A(counter[0]), .ZN(n_0_2));
   DFF_X1 finish_reg (.D(n_0_60), .CK(n_0_1), .Q(finish), .QN());
   DFF_X1 \A_reg[14]  (.D(n_0_20), .CK(n_0_1), .Q(A[14]), .QN());
   DFF_X1 \A_reg[13]  (.D(n_0_19), .CK(n_0_1), .Q(A[13]), .QN());
   DFF_X1 \A_reg[12]  (.D(n_0_18), .CK(n_0_1), .Q(A[12]), .QN());
   DFF_X1 \A_reg[11]  (.D(n_0_17), .CK(n_0_1), .Q(A[11]), .QN());
   DFF_X1 \A_reg[10]  (.D(n_0_16), .CK(n_0_1), .Q(A[10]), .QN());
   DFF_X1 \A_reg[9]  (.D(n_0_15), .CK(n_0_1), .Q(A[9]), .QN());
   DFF_X1 \A_reg[8]  (.D(n_0_14), .CK(n_0_1), .Q(A[8]), .QN());
   DFF_X1 \A_reg[7]  (.D(n_0_13), .CK(n_0_1), .Q(A[7]), .QN());
   DFF_X1 \A_reg[6]  (.D(n_0_12), .CK(n_0_1), .Q(A[6]), .QN());
   DFF_X1 \A_reg[5]  (.D(n_0_11), .CK(n_0_1), .Q(A[5]), .QN());
   DFF_X1 \A_reg[4]  (.D(n_0_10), .CK(n_0_1), .Q(A[4]), .QN());
   DFF_X1 \A_reg[3]  (.D(n_0_9), .CK(n_0_1), .Q(A[3]), .QN());
   DFF_X1 \A_reg[2]  (.D(n_0_8), .CK(n_0_1), .Q(A[2]), .QN());
   DFF_X1 \A_reg[1]  (.D(n_0_7), .CK(n_0_1), .Q(A[1]), .QN());
   DFF_X1 \A_reg[0]  (.D(n_0_6), .CK(n_0_1), .Q(A[0]), .QN());
   CLKGATETST_X1 clk_gate_multiplicand_buffer_reg (.CK(clk), .E(n_0_59), 
      .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \multiplicand_buffer_reg[15]  (.D(n_0_58), .CK(n_0_0), .Q(
      multiplicand_buffer[15]), .QN());
   DFF_X1 \multiplicand_buffer_reg[14]  (.D(n_0_57), .CK(n_0_0), .Q(
      multiplicand_buffer[14]), .QN());
   DFF_X1 \multiplicand_buffer_reg[13]  (.D(n_0_56), .CK(n_0_0), .Q(
      multiplicand_buffer[13]), .QN());
   DFF_X1 \multiplicand_buffer_reg[12]  (.D(n_0_55), .CK(n_0_0), .Q(
      multiplicand_buffer[12]), .QN());
   DFF_X1 \multiplicand_buffer_reg[11]  (.D(n_0_54), .CK(n_0_0), .Q(
      multiplicand_buffer[11]), .QN());
   DFF_X1 \multiplicand_buffer_reg[10]  (.D(n_0_53), .CK(n_0_0), .Q(
      multiplicand_buffer[10]), .QN());
   DFF_X1 \multiplicand_buffer_reg[9]  (.D(n_0_52), .CK(n_0_0), .Q(
      multiplicand_buffer[9]), .QN());
   DFF_X1 \multiplicand_buffer_reg[8]  (.D(n_0_51), .CK(n_0_0), .Q(
      multiplicand_buffer[8]), .QN());
   DFF_X1 \multiplicand_buffer_reg[7]  (.D(n_0_50), .CK(n_0_0), .Q(
      multiplicand_buffer[7]), .QN());
   DFF_X1 \multiplicand_buffer_reg[6]  (.D(n_0_49), .CK(n_0_0), .Q(
      multiplicand_buffer[6]), .QN());
   DFF_X1 \multiplicand_buffer_reg[5]  (.D(n_0_48), .CK(n_0_0), .Q(
      multiplicand_buffer[5]), .QN());
   DFF_X1 \multiplicand_buffer_reg[4]  (.D(n_0_47), .CK(n_0_0), .Q(
      multiplicand_buffer[4]), .QN());
   DFF_X1 \multiplicand_buffer_reg[3]  (.D(n_0_46), .CK(n_0_0), .Q(
      multiplicand_buffer[3]), .QN());
   DFF_X1 \multiplicand_buffer_reg[2]  (.D(n_0_45), .CK(n_0_0), .Q(
      multiplicand_buffer[2]), .QN());
   DFF_X1 \multiplicand_buffer_reg[1]  (.D(n_0_44), .CK(n_0_0), .Q(
      multiplicand_buffer[1]), .QN());
   DFF_X1 \multiplicand_buffer_reg[0]  (.D(n_0_43), .CK(n_0_0), .Q(
      multiplicand_buffer[0]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_0_37), .CK(n_0_1), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_0_36), .CK(n_0_1), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_0_35), .CK(n_0_1), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_0_34), .CK(n_0_1), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_0_33), .CK(n_0_1), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_0_32), .CK(n_0_1), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_0_31), .CK(n_0_1), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_0_30), .CK(n_0_1), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_0_29), .CK(n_0_1), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_0_28), .CK(n_0_1), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_0_27), .CK(n_0_1), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_0_26), .CK(n_0_1), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_0_25), .CK(n_0_1), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_0_24), .CK(n_0_1), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_0_23), .CK(n_0_1), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_0_22), .CK(n_0_1), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0_21), .CK(n_0_1), .Q(Q[0]), .QN());
   DFF_X1 \counter_reg[2]  (.D(n_0_41), .CK(n_0_1), .Q(counter[2]), .QN());
   DFF_X1 \counter_reg[1]  (.D(n_0_40), .CK(n_0_1), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(n_0_39), .CK(n_0_1), .Q(counter[0]), .QN());
   DFF_X1 working_reg (.D(n_0_38), .CK(n_0_1), .Q(working), .QN());
   DFF_X1 start_buffer_reg (.D(n_0_3), .CK(clk), .Q(start_buffer), .QN());
   MUX2_X1 start_buffer_reg_enable_mux_0 (.A(start_buffer), .B(n_0_4), .S(n_0_5), 
      .Z(n_0_3));
   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_0_42), .SE(1'b0), .GCK(n_0_1));
   AOI21_X1 i_0_0_0 (.A(n_0_0_0), .B1(n_0_0_1), .B2(n_0_0_81), .ZN(n_0_6));
   OAI21_X1 i_0_0_1 (.A(n_0_0_22), .B1(n_0_0_1), .B2(n_0_0_81), .ZN(n_0_0_0));
   NAND2_X1 i_0_0_2 (.A1(n_0_0_82), .A2(n_0_0_79), .ZN(n_0_0_1));
   AOI211_X1 i_0_0_3 (.A(n_0_59), .B(n_0_0_2), .C1(n_0_0_64), .C2(n_0_0_73), 
      .ZN(n_0_7));
   AOI22_X1 i_0_0_4 (.A1(n_0_0_80), .A2(n_0_0_79), .B1(n_0_0_75), .B2(n_0_0_73), 
      .ZN(n_0_0_2));
   AOI21_X1 i_0_0_5 (.A(n_0_0_3), .B1(n_0_0_31), .B2(n_0_0_72), .ZN(n_0_8));
   OAI21_X1 i_0_0_6 (.A(n_0_0_22), .B1(n_0_0_72), .B2(n_0_0_31), .ZN(n_0_0_3));
   AOI21_X1 i_0_0_7 (.A(n_0_0_5), .B1(n_0_0_50), .B2(n_0_0_71), .ZN(n_0_9));
   OAI21_X1 i_0_0_8 (.A(n_0_0_22), .B1(n_0_0_71), .B2(n_0_0_50), .ZN(n_0_0_5));
   AOI21_X1 i_0_0_9 (.A(n_0_0_7), .B1(n_0_0_8), .B2(n_0_0_84), .ZN(n_0_10));
   OAI21_X1 i_0_0_10 (.A(n_0_0_22), .B1(n_0_0_8), .B2(n_0_0_84), .ZN(n_0_0_7));
   XNOR2_X1 i_0_0_11 (.A(A[6]), .B(n_0_0_70), .ZN(n_0_0_8));
   AOI21_X1 i_0_0_12 (.A(n_0_0_91), .B1(n_0_0_96), .B2(n_0_0_92), .ZN(n_0_12));
   AOI21_X1 i_0_0_13 (.A(n_0_0_23), .B1(n_0_0_24), .B2(n_0_0_32), .ZN(n_0_18));
   OAI21_X1 i_0_0_14 (.A(n_0_0_22), .B1(n_0_0_32), .B2(n_0_0_24), .ZN(n_0_0_23));
   NAND2_X1 i_0_0_15 (.A1(n_0_0_28), .A2(n_0_0_27), .ZN(n_0_0_24));
   AOI21_X1 i_0_0_16 (.A(n_0_0_25), .B1(n_0_0_26), .B2(n_0_0_182), .ZN(n_0_19));
   OAI21_X1 i_0_0_17 (.A(n_0_0_22), .B1(n_0_0_182), .B2(n_0_0_26), .ZN(n_0_0_25));
   MUX2_X1 i_0_0_18 (.A(n_0_0_28), .B(n_0_0_27), .S(n_0_0_32), .Z(n_0_0_26));
   NAND2_X1 i_0_0_19 (.A1(n_0_0_15), .A2(n_0_0_173), .ZN(n_0_0_27));
   OR2_X1 i_0_0_20 (.A1(n_0_0_15), .A2(n_0_0_173), .ZN(n_0_0_28));
   AOI21_X1 i_0_0_21 (.A(n_0_0_140), .B1(n_0_0_167), .B2(n_0_0_141), .ZN(
      n_0_0_32));
   INV_X1 i_0_0_22 (.A(n_0_0_74), .ZN(n_0_0_64));
   AOI221_X1 i_0_0_23 (.A(n_0_0_69), .B1(n_0_0_41), .B2(multiplicand_buffer[2]), 
      .C1(multiplicand_buffer[3]), .C2(n_0_0_40), .ZN(n_0_0_17));
   NOR2_X1 i_0_0_24 (.A1(n_0_0_46), .A2(n_0_0_77), .ZN(n_0_0_69));
   OAI221_X1 i_0_0_25 (.A(n_0_0_76), .B1(n_0_0_46), .B2(n_0_0_176), .C1(n_0_0_38), 
      .C2(n_0_0_77), .ZN(n_0_0_18));
   NAND2_X1 i_0_0_26 (.A1(multiplicand_buffer[1]), .A2(n_0_0_41), .ZN(n_0_0_76));
   XOR2_X1 i_0_0_27 (.A(multiplicand_buffer[2]), .B(n_0_0_177), .Z(n_0_0_77));
   AOI21_X1 i_0_0_28 (.A(n_0_59), .B1(n_0_0_146), .B2(n_0_0_130), .ZN(n_0_20));
   OAI211_X1 i_0_0_29 (.A(n_0_0_131), .B(Q[2]), .C1(A[14]), .C2(n_0_0_42), 
      .ZN(n_0_0_130));
   NAND2_X1 i_0_0_30 (.A1(n_0_0_186), .A2(n_0_0_42), .ZN(n_0_0_131));
   OAI21_X1 i_0_0_31 (.A(n_0_0_147), .B1(n_0_0_48), .B2(multiplicand_buffer[15]), 
      .ZN(n_0_0_146));
   AOI21_X1 i_0_0_32 (.A(Q[2]), .B1(n_0_0_48), .B2(n_0_0_15), .ZN(n_0_0_147));
   AND2_X1 i_0_0_164 (.A1(Q[2]), .A2(n_0_0_22), .ZN(n_0_21));
   INV_X1 i_0_0_33 (.A(n_0_0_148), .ZN(n_0_22));
   AOI22_X1 i_0_0_34 (.A1(Q[3]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[0]), 
      .ZN(n_0_0_148));
   INV_X1 i_0_0_167 (.A(n_0_0_149), .ZN(n_0_23));
   AOI22_X1 i_0_0_168 (.A1(Q[4]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[1]), 
      .ZN(n_0_0_149));
   INV_X1 i_0_0_169 (.A(n_0_0_150), .ZN(n_0_24));
   AOI22_X1 i_0_0_170 (.A1(Q[5]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[2]), 
      .ZN(n_0_0_150));
   INV_X1 i_0_0_171 (.A(n_0_0_151), .ZN(n_0_25));
   AOI22_X1 i_0_0_172 (.A1(Q[6]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[3]), 
      .ZN(n_0_0_151));
   INV_X1 i_0_0_173 (.A(n_0_0_152), .ZN(n_0_26));
   AOI22_X1 i_0_0_174 (.A1(Q[7]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[4]), 
      .ZN(n_0_0_152));
   INV_X1 i_0_0_175 (.A(n_0_0_153), .ZN(n_0_27));
   AOI22_X1 i_0_0_176 (.A1(Q[8]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[5]), 
      .ZN(n_0_0_153));
   INV_X1 i_0_0_177 (.A(n_0_0_154), .ZN(n_0_28));
   AOI22_X1 i_0_0_178 (.A1(Q[9]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[6]), 
      .ZN(n_0_0_154));
   INV_X1 i_0_0_179 (.A(n_0_0_155), .ZN(n_0_29));
   AOI22_X1 i_0_0_180 (.A1(Q[10]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[7]), 
      .ZN(n_0_0_155));
   INV_X1 i_0_0_181 (.A(n_0_0_156), .ZN(n_0_30));
   AOI22_X1 i_0_0_182 (.A1(Q[11]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[8]), 
      .ZN(n_0_0_156));
   INV_X1 i_0_0_183 (.A(n_0_0_157), .ZN(n_0_31));
   AOI22_X1 i_0_0_184 (.A1(Q[12]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[9]), 
      .ZN(n_0_0_157));
   INV_X1 i_0_0_185 (.A(n_0_0_158), .ZN(n_0_32));
   AOI22_X1 i_0_0_186 (.A1(Q[13]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[10]), 
      .ZN(n_0_0_158));
   INV_X1 i_0_0_187 (.A(n_0_0_159), .ZN(n_0_33));
   AOI22_X1 i_0_0_188 (.A1(Q[14]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[11]), 
      .ZN(n_0_0_159));
   INV_X1 i_0_0_189 (.A(n_0_0_160), .ZN(n_0_34));
   AOI22_X1 i_0_0_190 (.A1(Q[15]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[12]), 
      .ZN(n_0_0_160));
   INV_X1 i_0_0_191 (.A(n_0_0_161), .ZN(n_0_35));
   AOI22_X1 i_0_0_192 (.A1(Q[16]), .A2(n_0_0_22), .B1(n_0_4), .B2(multiplier[13]), 
      .ZN(n_0_0_161));
   INV_X1 i_0_0_35 (.A(n_0_0_162), .ZN(n_0_36));
   AOI22_X1 i_0_0_36 (.A1(n_0_0_163), .A2(n_0_0_164), .B1(n_0_4), .B2(
      multiplier[14]), .ZN(n_0_0_162));
   NOR2_X1 i_0_0_37 (.A1(n_0_0_179), .A2(n_0_59), .ZN(n_0_0_163));
   NAND2_X1 i_0_0_38 (.A1(n_0_0_14), .A2(n_0_0_180), .ZN(n_0_0_164));
   INV_X1 i_0_0_39 (.A(n_0_0_165), .ZN(n_0_37));
   AOI22_X1 i_0_0_40 (.A1(n_0_0_166), .A2(n_0_0_19), .B1(n_0_4), .B2(
      multiplier[15]), .ZN(n_0_0_165));
   NOR2_X1 i_0_0_41 (.A1(n_0_0_168), .A2(n_0_59), .ZN(n_0_0_166));
   NAND2_X1 i_0_0_42 (.A1(n_0_0_179), .A2(n_0_0_169), .ZN(n_0_0_19));
   NOR2_X1 i_0_0_43 (.A1(n_0_0_179), .A2(n_0_0_169), .ZN(n_0_0_168));
   XNOR2_X1 i_0_0_44 (.A(A[1]), .B(n_0_0_20), .ZN(n_0_0_169));
   AOI221_X1 i_0_0_45 (.A(n_0_0_175), .B1(n_0_0_40), .B2(multiplicand_buffer[1]), 
      .C1(n_0_0_171), .C2(multiplicand_buffer[0]), .ZN(n_0_0_20));
   OAI21_X1 i_0_0_46 (.A(n_0_0_46), .B1(n_0_0_42), .B2(Q[2]), .ZN(n_0_0_171));
   NOR2_X1 i_0_0_47 (.A1(n_0_0_38), .A2(n_0_0_176), .ZN(n_0_0_175));
   XNOR2_X1 i_0_0_48 (.A(multiplicand_buffer[1]), .B(multiplicand_buffer[0]), 
      .ZN(n_0_0_176));
   NOR2_X1 i_0_0_49 (.A1(multiplicand_buffer[1]), .A2(multiplicand_buffer[0]), 
      .ZN(n_0_0_177));
   NOR2_X1 i_0_0_50 (.A1(n_0_0_14), .A2(n_0_0_180), .ZN(n_0_0_179));
   NAND3_X1 i_0_0_51 (.A1(n_0_0_47), .A2(multiplicand_buffer[0]), .A3(n_0_0_42), 
      .ZN(n_0_0_180));
   AOI21_X1 i_0_0_52 (.A(rst), .B1(n_0_0_188), .B2(n_0_0_16), .ZN(n_0_38));
   NOR2_X1 i_0_0_53 (.A1(n_0_0_16), .A2(rst), .ZN(n_0_4));
   AND2_X1 i_0_0_219 (.A1(n_0_2), .A2(n_0_0_22), .ZN(n_0_39));
   AOI21_X1 i_0_0_54 (.A(n_0_0_184), .B1(counter[0]), .B2(counter[1]), .ZN(
      n_0_40));
   OAI21_X1 i_0_0_55 (.A(n_0_0_22), .B1(counter[0]), .B2(counter[1]), .ZN(
      n_0_0_184));
   NOR3_X1 i_0_0_56 (.A1(n_0_59), .A2(n_0_0_185), .A3(n_0_0_188), .ZN(n_0_41));
   AOI21_X1 i_0_0_57 (.A(counter[2]), .B1(counter[1]), .B2(counter[0]), .ZN(
      n_0_0_185));
   OR2_X1 i_0_0_224 (.A1(n_0_59), .A2(working), .ZN(n_0_42));
   NOR2_X1 i_0_0_58 (.A1(n_0_0_216), .A2(rst), .ZN(n_0_43));
   NOR2_X1 i_0_0_226 (.A1(n_0_0_217), .A2(rst), .ZN(n_0_44));
   NOR2_X1 i_0_0_227 (.A1(n_0_0_218), .A2(rst), .ZN(n_0_45));
   NOR2_X1 i_0_0_228 (.A1(n_0_0_219), .A2(rst), .ZN(n_0_46));
   NOR2_X1 i_0_0_229 (.A1(n_0_0_220), .A2(rst), .ZN(n_0_47));
   NOR2_X1 i_0_0_230 (.A1(n_0_0_221), .A2(rst), .ZN(n_0_48));
   NOR2_X1 i_0_0_231 (.A1(n_0_0_222), .A2(rst), .ZN(n_0_49));
   NOR2_X1 i_0_0_232 (.A1(n_0_0_223), .A2(rst), .ZN(n_0_50));
   NOR2_X1 i_0_0_233 (.A1(n_0_0_224), .A2(rst), .ZN(n_0_51));
   NOR2_X1 i_0_0_234 (.A1(n_0_0_225), .A2(rst), .ZN(n_0_52));
   NOR2_X1 i_0_0_235 (.A1(n_0_0_4), .A2(rst), .ZN(n_0_53));
   NOR2_X1 i_0_0_236 (.A1(n_0_0_6), .A2(rst), .ZN(n_0_54));
   NOR2_X1 i_0_0_237 (.A1(n_0_0_9), .A2(rst), .ZN(n_0_55));
   NOR2_X1 i_0_0_238 (.A1(n_0_0_10), .A2(rst), .ZN(n_0_56));
   NOR2_X1 i_0_0_239 (.A1(n_0_0_11), .A2(rst), .ZN(n_0_57));
   NOR2_X1 i_0_0_240 (.A1(n_0_0_12), .A2(rst), .ZN(n_0_58));
   AND2_X1 i_0_0_241 (.A1(n_0_0_188), .A2(n_0_0_22), .ZN(n_0_60));
   AND3_X1 i_0_0_59 (.A1(counter[2]), .A2(counter[1]), .A3(counter[0]), .ZN(
      n_0_0_188));
   AOI211_X1 i_0_0_246 (.A(n_0_0_13), .B(n_0_0_189), .C1(n_0_0_193), .C2(
      n_0_0_195), .ZN(overflow_flag));
   NOR4_X1 i_0_0_247 (.A1(n_0_0_15), .A2(n_0_0_192), .A3(n_0_0_191), .A4(
      n_0_0_190), .ZN(n_0_0_189));
   OAI211_X1 i_0_0_248 (.A(A[8]), .B(A[7]), .C1(A[6]), .C2(n_0_0_202), .ZN(
      n_0_0_190));
   NAND3_X1 i_0_0_249 (.A1(A[12]), .A2(A[10]), .A3(A[9]), .ZN(n_0_0_191));
   NAND2_X1 i_0_0_250 (.A1(A[13]), .A2(A[11]), .ZN(n_0_0_192));
   NOR4_X1 i_0_0_251 (.A1(n_0_0_194), .A2(A[9]), .A3(A[11]), .A4(A[14]), 
      .ZN(n_0_0_193));
   OR3_X1 i_0_0_252 (.A1(A[13]), .A2(A[12]), .A3(A[10]), .ZN(n_0_0_194));
   NOR4_X1 i_0_0_253 (.A1(A[8]), .A2(A[7]), .A3(A[6]), .A4(n_0_0_202), .ZN(
      n_0_0_195));
   XOR2_X1 i_0_0_254 (.A(Q[8]), .B(Q[7]), .Z(result[0]));
   NOR2_X1 i_0_0_60 (.A1(n_0_0_214), .A2(n_0_0_196), .ZN(result[1]));
   AOI21_X1 i_0_0_61 (.A(Q[9]), .B1(Q[8]), .B2(Q[7]), .ZN(n_0_0_196));
   XNOR2_X1 i_0_0_62 (.A(Q[10]), .B(n_0_0_215), .ZN(result[2]));
   XNOR2_X1 i_0_0_63 (.A(Q[11]), .B(n_0_0_213), .ZN(result[3]));
   NOR2_X1 i_0_0_64 (.A1(n_0_0_211), .A2(n_0_0_197), .ZN(result[4]));
   NOR2_X1 i_0_0_65 (.A1(Q[12]), .A2(n_0_0_212), .ZN(n_0_0_197));
   XOR2_X1 i_0_0_66 (.A(Q[13]), .B(n_0_0_211), .Z(result[5]));
   NOR2_X1 i_0_0_67 (.A1(n_0_0_210), .A2(n_0_0_198), .ZN(result[6]));
   AOI21_X1 i_0_0_68 (.A(Q[14]), .B1(Q[13]), .B2(n_0_0_211), .ZN(n_0_0_198));
   XOR2_X1 i_0_0_69 (.A(Q[15]), .B(n_0_0_210), .Z(result[7]));
   NOR2_X1 i_0_0_265 (.A1(n_0_0_208), .A2(n_0_0_199), .ZN(result[8]));
   AOI21_X1 i_0_0_266 (.A(Q[16]), .B1(Q[15]), .B2(n_0_0_210), .ZN(n_0_0_199));
   XNOR2_X1 i_0_0_267 (.A(A[0]), .B(n_0_0_209), .ZN(result[9]));
   XNOR2_X1 i_0_0_268 (.A(n_0_0_21), .B(n_0_0_207), .ZN(result[10]));
   NOR2_X1 i_0_0_269 (.A1(n_0_0_205), .A2(n_0_0_200), .ZN(result[11]));
   AOI21_X1 i_0_0_270 (.A(A[2]), .B1(A[1]), .B2(n_0_0_207), .ZN(n_0_0_200));
   XNOR2_X1 i_0_0_271 (.A(A[3]), .B(n_0_0_206), .ZN(result[12]));
   XOR2_X1 i_0_0_272 (.A(A[4]), .B(n_0_0_204), .Z(result[13]));
   NOR2_X1 i_0_0_273 (.A1(n_0_0_202), .A2(n_0_0_201), .ZN(result[14]));
   AOI21_X1 i_0_0_274 (.A(A[5]), .B1(A[4]), .B2(n_0_0_204), .ZN(n_0_0_201));
   XNOR2_X1 i_0_0_275 (.A(A[6]), .B(n_0_0_203), .ZN(result[15]));
   INV_X1 i_0_0_276 (.A(n_0_0_203), .ZN(n_0_0_202));
   NAND3_X1 i_0_0_277 (.A1(A[5]), .A2(A[4]), .A3(n_0_0_204), .ZN(n_0_0_203));
   AND2_X1 i_0_0_278 (.A1(A[3]), .A2(n_0_0_205), .ZN(n_0_0_204));
   INV_X1 i_0_0_279 (.A(n_0_0_206), .ZN(n_0_0_205));
   NAND3_X1 i_0_0_280 (.A1(A[2]), .A2(A[1]), .A3(n_0_0_207), .ZN(n_0_0_206));
   NOR2_X1 i_0_0_281 (.A1(n_0_0_14), .A2(n_0_0_209), .ZN(n_0_0_207));
   INV_X1 i_0_0_282 (.A(n_0_0_209), .ZN(n_0_0_208));
   NAND3_X1 i_0_0_283 (.A1(Q[16]), .A2(Q[15]), .A3(n_0_0_210), .ZN(n_0_0_209));
   AND3_X1 i_0_0_70 (.A1(Q[14]), .A2(Q[13]), .A3(n_0_0_211), .ZN(n_0_0_210));
   AND2_X1 i_0_0_71 (.A1(Q[12]), .A2(n_0_0_212), .ZN(n_0_0_211));
   AND3_X1 i_0_0_72 (.A1(Q[11]), .A2(Q[10]), .A3(n_0_0_214), .ZN(n_0_0_212));
   NAND2_X1 i_0_0_73 (.A1(Q[10]), .A2(n_0_0_214), .ZN(n_0_0_213));
   INV_X1 i_0_0_74 (.A(n_0_0_215), .ZN(n_0_0_214));
   NAND3_X1 i_0_0_75 (.A1(Q[9]), .A2(Q[8]), .A3(Q[7]), .ZN(n_0_0_215));
   INV_X1 i_0_0_76 (.A(multiplicand[0]), .ZN(n_0_0_216));
   INV_X1 i_0_0_291 (.A(multiplicand[1]), .ZN(n_0_0_217));
   INV_X1 i_0_0_292 (.A(multiplicand[2]), .ZN(n_0_0_218));
   INV_X1 i_0_0_293 (.A(multiplicand[3]), .ZN(n_0_0_219));
   INV_X1 i_0_0_294 (.A(multiplicand[4]), .ZN(n_0_0_220));
   INV_X1 i_0_0_295 (.A(multiplicand[5]), .ZN(n_0_0_221));
   INV_X1 i_0_0_296 (.A(multiplicand[6]), .ZN(n_0_0_222));
   INV_X1 i_0_0_297 (.A(multiplicand[7]), .ZN(n_0_0_223));
   INV_X1 i_0_0_298 (.A(multiplicand[8]), .ZN(n_0_0_224));
   INV_X1 i_0_0_299 (.A(multiplicand[9]), .ZN(n_0_0_225));
   INV_X1 i_0_0_300 (.A(multiplicand[10]), .ZN(n_0_0_4));
   INV_X1 i_0_0_301 (.A(multiplicand[11]), .ZN(n_0_0_6));
   INV_X1 i_0_0_302 (.A(multiplicand[12]), .ZN(n_0_0_9));
   INV_X1 i_0_0_303 (.A(multiplicand[13]), .ZN(n_0_0_10));
   INV_X1 i_0_0_304 (.A(multiplicand[14]), .ZN(n_0_0_11));
   INV_X1 i_0_0_305 (.A(multiplicand[15]), .ZN(n_0_0_12));
   INV_X1 i_0_0_307 (.A(finish), .ZN(n_0_0_13));
   INV_X1 i_0_0_77 (.A(A[0]), .ZN(n_0_0_14));
   INV_X1 i_0_0_78 (.A(A[1]), .ZN(n_0_0_21));
   INV_X1 i_0_0_79 (.A(A[14]), .ZN(n_0_0_15));
   INV_X1 i_0_0_80 (.A(n_0_0_29), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_81 (.A1(start), .A2(n_0_0_22), .ZN(n_0_5));
   NOR2_X1 i_0_0_82 (.A1(rst), .A2(n_0_0_29), .ZN(n_0_0_22));
   NOR2_X1 i_0_0_83 (.A1(start_buffer), .A2(n_0_0_30), .ZN(n_0_0_29));
   INV_X1 i_0_0_84 (.A(start), .ZN(n_0_0_30));
   AOI21_X1 i_0_0_85 (.A(n_0_0_34), .B1(A[4]), .B2(n_0_0_36), .ZN(n_0_0_31));
   INV_X1 i_0_0_86 (.A(n_0_0_34), .ZN(n_0_0_33));
   NOR2_X1 i_0_0_87 (.A1(A[4]), .A2(n_0_0_36), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_88 (.A1(A[4]), .A2(n_0_0_36), .ZN(n_0_0_35));
   OAI221_X1 i_0_0_89 (.A(n_0_0_37), .B1(n_0_0_46), .B2(n_0_0_43), .C1(n_0_0_39), 
      .C2(n_0_0_38), .ZN(n_0_0_36));
   AOI22_X1 i_0_0_90 (.A1(multiplicand_buffer[4]), .A2(n_0_0_40), .B1(
      multiplicand_buffer[3]), .B2(n_0_0_41), .ZN(n_0_0_37));
   NAND3_X1 i_0_0_91 (.A1(Q[2]), .A2(n_0_0_42), .A3(n_0_0_47), .ZN(n_0_0_38));
   XNOR2_X1 i_0_0_92 (.A(multiplicand_buffer[4]), .B(n_0_0_44), .ZN(n_0_0_39));
   AOI211_X1 i_0_0_93 (.A(Q[2]), .B(n_0_0_48), .C1(Q[1]), .C2(Q[0]), .ZN(
      n_0_0_40));
   NOR2_X1 i_0_0_94 (.A1(Q[2]), .A2(n_0_0_42), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_95 (.A1(Q[1]), .A2(Q[0]), .ZN(n_0_0_42));
   OAI21_X1 i_0_0_96 (.A(n_0_0_44), .B1(n_0_0_49), .B2(n_0_0_45), .ZN(n_0_0_43));
   NAND2_X1 i_0_0_97 (.A1(n_0_0_49), .A2(n_0_0_45), .ZN(n_0_0_44));
   NOR3_X1 i_0_0_98 (.A1(multiplicand_buffer[2]), .A2(multiplicand_buffer[0]), 
      .A3(multiplicand_buffer[1]), .ZN(n_0_0_45));
   NAND2_X1 i_0_0_99 (.A1(Q[2]), .A2(n_0_0_48), .ZN(n_0_0_46));
   INV_X1 i_0_0_100 (.A(n_0_0_48), .ZN(n_0_0_47));
   NOR2_X1 i_0_0_101 (.A1(Q[1]), .A2(Q[0]), .ZN(n_0_0_48));
   INV_X1 i_0_0_102 (.A(multiplicand_buffer[3]), .ZN(n_0_0_49));
   OAI21_X1 i_0_0_103 (.A(n_0_0_52), .B1(A[5]), .B2(n_0_0_53), .ZN(n_0_0_50));
   NOR2_X1 i_0_0_104 (.A1(A[5]), .A2(n_0_0_53), .ZN(n_0_0_51));
   NAND2_X1 i_0_0_105 (.A1(A[5]), .A2(n_0_0_53), .ZN(n_0_0_52));
   OAI221_X1 i_0_0_106 (.A(n_0_0_54), .B1(n_0_0_46), .B2(n_0_0_39), .C1(n_0_0_38), 
      .C2(n_0_0_55), .ZN(n_0_0_53));
   AOI22_X1 i_0_0_107 (.A1(multiplicand_buffer[5]), .A2(n_0_0_40), .B1(n_0_0_41), 
      .B2(multiplicand_buffer[4]), .ZN(n_0_0_54));
   XOR2_X1 i_0_0_108 (.A(multiplicand_buffer[5]), .B(n_0_0_56), .Z(n_0_0_55));
   NOR2_X1 i_0_0_109 (.A1(multiplicand_buffer[4]), .A2(n_0_0_44), .ZN(n_0_0_56));
   INV_X1 i_0_0_110 (.A(multiplicand_buffer[5]), .ZN(n_0_0_57));
   AOI21_X1 i_0_0_111 (.A(n_0_0_58), .B1(n_0_0_66), .B2(n_0_0_59), .ZN(n_0_11));
   OAI21_X1 i_0_0_112 (.A(n_0_0_22), .B1(n_0_0_66), .B2(n_0_0_59), .ZN(n_0_0_58));
   OAI21_X1 i_0_0_113 (.A(n_0_0_61), .B1(A[7]), .B2(n_0_0_62), .ZN(n_0_0_59));
   NOR2_X1 i_0_0_114 (.A1(A[7]), .A2(n_0_0_62), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_115 (.A1(A[7]), .A2(n_0_0_62), .ZN(n_0_0_61));
   OAI221_X1 i_0_0_116 (.A(n_0_0_63), .B1(n_0_0_46), .B2(n_0_0_86), .C1(n_0_0_38), 
      .C2(n_0_0_65), .ZN(n_0_0_62));
   AOI22_X1 i_0_0_117 (.A1(multiplicand_buffer[7]), .A2(n_0_0_40), .B1(
      multiplicand_buffer[6]), .B2(n_0_0_41), .ZN(n_0_0_63));
   XOR2_X1 i_0_0_118 (.A(multiplicand_buffer[7]), .B(n_0_0_88), .Z(n_0_0_65));
   OAI21_X1 i_0_0_119 (.A(n_0_0_67), .B1(A[6]), .B2(n_0_0_70), .ZN(n_0_0_66));
   NAND2_X1 i_0_0_120 (.A1(n_0_0_84), .A2(n_0_0_68), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_121 (.A1(A[6]), .A2(n_0_0_70), .ZN(n_0_0_68));
   AOI21_X1 i_0_0_122 (.A(n_0_0_51), .B1(n_0_0_52), .B2(n_0_0_71), .ZN(n_0_0_70));
   OAI21_X1 i_0_0_123 (.A(n_0_0_33), .B1(n_0_0_90), .B2(n_0_0_72), .ZN(n_0_0_71));
   NAND2_X1 i_0_0_124 (.A1(n_0_0_74), .A2(n_0_0_73), .ZN(n_0_0_72));
   NAND2_X1 i_0_0_125 (.A1(A[3]), .A2(n_0_0_78), .ZN(n_0_0_73));
   NAND3_X1 i_0_0_126 (.A1(n_0_0_80), .A2(n_0_0_79), .A3(n_0_0_75), .ZN(n_0_0_74));
   OR2_X1 i_0_0_127 (.A1(A[3]), .A2(n_0_0_78), .ZN(n_0_0_75));
   OAI21_X1 i_0_0_128 (.A(n_0_0_17), .B1(n_0_0_38), .B2(n_0_0_43), .ZN(n_0_0_78));
   OR2_X1 i_0_0_129 (.A1(A[2]), .A2(n_0_0_83), .ZN(n_0_0_79));
   NAND2_X1 i_0_0_130 (.A1(n_0_0_82), .A2(n_0_0_81), .ZN(n_0_0_80));
   AOI21_X1 i_0_0_131 (.A(n_0_0_18), .B1(multiplicand_buffer[2]), .B2(n_0_0_40), 
      .ZN(n_0_0_81));
   NAND2_X1 i_0_0_132 (.A1(A[2]), .A2(n_0_0_83), .ZN(n_0_0_82));
   OAI21_X1 i_0_0_133 (.A(n_0_0_19), .B1(n_0_0_20), .B2(n_0_0_21), .ZN(n_0_0_83));
   AOI221_X1 i_0_0_134 (.A(n_0_0_85), .B1(multiplicand_buffer[5]), .B2(n_0_0_41), 
      .C1(multiplicand_buffer[6]), .C2(n_0_0_40), .ZN(n_0_0_84));
   OAI22_X1 i_0_0_135 (.A1(n_0_0_38), .A2(n_0_0_86), .B1(n_0_0_55), .B2(n_0_0_46), 
      .ZN(n_0_0_85));
   INV_X1 i_0_0_136 (.A(n_0_0_87), .ZN(n_0_0_86));
   AOI21_X1 i_0_0_137 (.A(n_0_0_88), .B1(multiplicand_buffer[6]), .B2(n_0_0_89), 
      .ZN(n_0_0_87));
   NOR2_X1 i_0_0_138 (.A1(multiplicand_buffer[6]), .A2(n_0_0_89), .ZN(n_0_0_88));
   NAND2_X1 i_0_0_139 (.A1(n_0_0_56), .A2(n_0_0_57), .ZN(n_0_0_89));
   INV_X1 i_0_0_140 (.A(n_0_0_35), .ZN(n_0_0_90));
   OAI21_X1 i_0_0_141 (.A(n_0_0_22), .B1(n_0_0_96), .B2(n_0_0_92), .ZN(n_0_0_91));
   OAI221_X1 i_0_0_142 (.A(n_0_0_93), .B1(n_0_0_46), .B2(n_0_0_65), .C1(n_0_0_38), 
      .C2(n_0_0_94), .ZN(n_0_0_92));
   AOI22_X1 i_0_0_143 (.A1(n_0_0_41), .A2(multiplicand_buffer[7]), .B1(
      multiplicand_buffer[8]), .B2(n_0_0_40), .ZN(n_0_0_93));
   XOR2_X1 i_0_0_144 (.A(multiplicand_buffer[8]), .B(n_0_0_95), .Z(n_0_0_94));
   NOR3_X1 i_0_0_145 (.A1(multiplicand_buffer[6]), .A2(n_0_0_89), .A3(
      multiplicand_buffer[7]), .ZN(n_0_0_95));
   XOR2_X1 i_0_0_146 (.A(A[8]), .B(n_0_0_97), .Z(n_0_0_96));
   AOI21_X1 i_0_0_147 (.A(n_0_0_60), .B1(n_0_0_66), .B2(n_0_0_61), .ZN(n_0_0_97));
   INV_X1 i_0_0_148 (.A(multiplicand_buffer[8]), .ZN(n_0_0_98));
   AOI21_X1 i_0_0_149 (.A(n_0_0_99), .B1(n_0_0_108), .B2(n_0_0_100), .ZN(n_0_13));
   OAI21_X1 i_0_0_150 (.A(n_0_0_22), .B1(n_0_0_108), .B2(n_0_0_100), .ZN(
      n_0_0_99));
   NAND2_X1 i_0_0_151 (.A1(n_0_0_102), .A2(n_0_0_101), .ZN(n_0_0_100));
   OR2_X1 i_0_0_152 (.A1(A[9]), .A2(n_0_0_103), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_153 (.A1(A[9]), .A2(n_0_0_103), .ZN(n_0_0_102));
   OAI221_X1 i_0_0_154 (.A(n_0_0_104), .B1(n_0_0_94), .B2(n_0_0_46), .C1(
      n_0_0_38), .C2(n_0_0_105), .ZN(n_0_0_103));
   AOI22_X1 i_0_0_155 (.A1(multiplicand_buffer[9]), .A2(n_0_0_40), .B1(
      multiplicand_buffer[8]), .B2(n_0_0_41), .ZN(n_0_0_104));
   OAI21_X1 i_0_0_156 (.A(n_0_0_106), .B1(n_0_0_110), .B2(n_0_0_107), .ZN(
      n_0_0_105));
   NAND2_X1 i_0_0_157 (.A1(n_0_0_110), .A2(n_0_0_107), .ZN(n_0_0_106));
   AND2_X1 i_0_0_158 (.A1(n_0_0_95), .A2(n_0_0_98), .ZN(n_0_0_107));
   AOI22_X1 i_0_0_159 (.A1(n_0_0_92), .A2(A[8]), .B1(n_0_0_97), .B2(n_0_0_109), 
      .ZN(n_0_0_108));
   OR2_X1 i_0_0_160 (.A1(n_0_0_92), .A2(A[8]), .ZN(n_0_0_109));
   INV_X1 i_0_0_161 (.A(multiplicand_buffer[9]), .ZN(n_0_0_110));
   AOI21_X1 i_0_0_162 (.A(n_0_0_111), .B1(n_0_0_118), .B2(n_0_0_112), .ZN(n_0_14));
   OAI21_X1 i_0_0_163 (.A(n_0_0_22), .B1(n_0_0_118), .B2(n_0_0_112), .ZN(
      n_0_0_111));
   OAI21_X1 i_0_0_165 (.A(n_0_0_114), .B1(A[10]), .B2(n_0_0_115), .ZN(n_0_0_112));
   NOR2_X1 i_0_0_166 (.A1(A[10]), .A2(n_0_0_115), .ZN(n_0_0_113));
   NAND2_X1 i_0_0_193 (.A1(A[10]), .A2(n_0_0_115), .ZN(n_0_0_114));
   OAI221_X1 i_0_0_194 (.A(n_0_0_116), .B1(n_0_0_46), .B2(n_0_0_105), .C1(
      n_0_0_38), .C2(n_0_0_117), .ZN(n_0_0_115));
   AOI22_X1 i_0_0_195 (.A1(n_0_0_41), .A2(multiplicand_buffer[9]), .B1(
      multiplicand_buffer[10]), .B2(n_0_0_40), .ZN(n_0_0_116));
   XNOR2_X1 i_0_0_196 (.A(multiplicand_buffer[10]), .B(n_0_0_106), .ZN(n_0_0_117));
   NAND2_X1 i_0_0_197 (.A1(n_0_0_101), .A2(n_0_0_119), .ZN(n_0_0_118));
   NAND2_X1 i_0_0_198 (.A1(n_0_0_102), .A2(n_0_0_108), .ZN(n_0_0_119));
   AOI211_X1 i_0_0_199 (.A(n_0_0_120), .B(n_0_59), .C1(n_0_0_126), .C2(n_0_0_121), 
      .ZN(n_0_15));
   NOR2_X1 i_0_0_200 (.A1(n_0_0_126), .A2(n_0_0_121), .ZN(n_0_0_120));
   XOR2_X1 i_0_0_201 (.A(A[11]), .B(n_0_0_122), .Z(n_0_0_121));
   OAI221_X1 i_0_0_202 (.A(n_0_0_123), .B1(n_0_0_46), .B2(n_0_0_117), .C1(
      n_0_0_38), .C2(n_0_0_124), .ZN(n_0_0_122));
   AOI22_X1 i_0_0_203 (.A1(n_0_0_41), .A2(multiplicand_buffer[10]), .B1(
      multiplicand_buffer[11]), .B2(n_0_0_40), .ZN(n_0_0_123));
   XOR2_X1 i_0_0_204 (.A(multiplicand_buffer[11]), .B(n_0_0_125), .Z(n_0_0_124));
   NOR2_X1 i_0_0_205 (.A1(multiplicand_buffer[10]), .A2(n_0_0_106), .ZN(
      n_0_0_125));
   AOI21_X1 i_0_0_206 (.A(n_0_0_113), .B1(n_0_0_118), .B2(n_0_0_114), .ZN(
      n_0_0_126));
   INV_X1 i_0_0_207 (.A(n_0_0_22), .ZN(n_0_59));
   NOR3_X1 i_0_0_208 (.A1(multiplicand_buffer[10]), .A2(n_0_0_106), .A3(
      multiplicand_buffer[11]), .ZN(n_0_0_127));
   XOR2_X1 i_0_0_209 (.A(multiplicand_buffer[12]), .B(n_0_0_127), .Z(n_0_0_128));
   AOI22_X1 i_0_0_210 (.A1(n_0_0_41), .A2(multiplicand_buffer[11]), .B1(n_0_0_40), 
      .B2(multiplicand_buffer[12]), .ZN(n_0_0_129));
   OAI221_X1 i_0_0_211 (.A(n_0_0_129), .B1(n_0_0_46), .B2(n_0_0_124), .C1(
      n_0_0_128), .C2(n_0_0_38), .ZN(n_0_0_132));
   OR2_X1 i_0_0_212 (.A1(n_0_0_122), .A2(A[11]), .ZN(n_0_0_133));
   AOI22_X1 i_0_0_213 (.A1(n_0_0_133), .A2(n_0_0_126), .B1(n_0_0_122), .B2(A[11]), 
      .ZN(n_0_0_134));
   XNOR2_X1 i_0_0_214 (.A(n_0_0_134), .B(A[12]), .ZN(n_0_0_135));
   OAI21_X1 i_0_0_215 (.A(n_0_0_22), .B1(n_0_0_132), .B2(n_0_0_135), .ZN(
      n_0_0_136));
   AOI21_X1 i_0_0_216 (.A(n_0_0_136), .B1(n_0_0_132), .B2(n_0_0_135), .ZN(n_0_16));
   INV_X1 i_0_0_217 (.A(multiplicand_buffer[12]), .ZN(n_0_0_137));
   AOI21_X1 i_0_0_218 (.A(n_0_0_138), .B1(n_0_0_167), .B2(n_0_0_139), .ZN(n_0_17));
   OAI21_X1 i_0_0_220 (.A(n_0_0_22), .B1(n_0_0_167), .B2(n_0_0_139), .ZN(
      n_0_0_138));
   OAI21_X1 i_0_0_221 (.A(n_0_0_141), .B1(A[13]), .B2(n_0_0_142), .ZN(n_0_0_139));
   NOR2_X1 i_0_0_222 (.A1(A[13]), .A2(n_0_0_142), .ZN(n_0_0_140));
   NAND2_X1 i_0_0_223 (.A1(A[13]), .A2(n_0_0_142), .ZN(n_0_0_141));
   OAI221_X1 i_0_0_225 (.A(n_0_0_143), .B1(n_0_0_128), .B2(n_0_0_46), .C1(
      n_0_0_38), .C2(n_0_0_144), .ZN(n_0_0_142));
   AOI22_X1 i_0_0_242 (.A1(multiplicand_buffer[13]), .A2(n_0_0_40), .B1(
      multiplicand_buffer[12]), .B2(n_0_0_41), .ZN(n_0_0_143));
   XNOR2_X1 i_0_0_243 (.A(multiplicand_buffer[13]), .B(n_0_0_145), .ZN(n_0_0_144));
   NAND2_X1 i_0_0_244 (.A1(n_0_0_127), .A2(n_0_0_137), .ZN(n_0_0_145));
   OAI21_X1 i_0_0_245 (.A(n_0_0_170), .B1(A[12]), .B2(n_0_0_132), .ZN(n_0_0_167));
   NAND2_X1 i_0_0_255 (.A1(n_0_0_134), .A2(n_0_0_172), .ZN(n_0_0_170));
   NAND2_X1 i_0_0_256 (.A1(A[12]), .A2(n_0_0_132), .ZN(n_0_0_172));
   OAI221_X1 i_0_0_257 (.A(n_0_0_174), .B1(n_0_0_46), .B2(n_0_0_144), .C1(
      n_0_0_38), .C2(n_0_0_178), .ZN(n_0_0_173));
   AOI22_X1 i_0_0_258 (.A1(multiplicand_buffer[14]), .A2(n_0_0_40), .B1(n_0_0_41), 
      .B2(multiplicand_buffer[13]), .ZN(n_0_0_174));
   XOR2_X1 i_0_0_259 (.A(multiplicand_buffer[14]), .B(n_0_0_181), .Z(n_0_0_178));
   NOR2_X1 i_0_0_260 (.A1(multiplicand_buffer[13]), .A2(n_0_0_145), .ZN(
      n_0_0_181));
   AOI221_X1 i_0_0_261 (.A(n_0_0_183), .B1(multiplicand_buffer[15]), .B2(
      n_0_0_40), .C1(multiplicand_buffer[14]), .C2(n_0_0_41), .ZN(n_0_0_182));
   OAI22_X1 i_0_0_262 (.A1(n_0_0_38), .A2(n_0_0_186), .B1(n_0_0_178), .B2(
      n_0_0_46), .ZN(n_0_0_183));
   XOR2_X1 i_0_0_263 (.A(multiplicand_buffer[15]), .B(n_0_0_187), .Z(n_0_0_186));
   NOR3_X1 i_0_0_264 (.A1(multiplicand_buffer[13]), .A2(n_0_0_145), .A3(
      multiplicand_buffer[14]), .ZN(n_0_0_187));
endmodule
