/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Apr 23 16:48:56 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1841939902 */

module adder(A, B, is_subtract, result, carry, overflow_flag, negative);
   input [15:0]A;
   input [15:0]B;
   input is_subtract;
   output [15:0]result;
   output carry;
   output overflow_flag;
   output negative;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_37;
   wire n_0_0_42;
   wire n_0_0_46;
   wire n_0_0_50;
   wire n_0_0_53;
   wire n_0_0_55;
   wire n_0_0_58;
   wire n_0_0_63;
   wire n_0_0_68;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_23;
   wire n_0_0_43;
   wire n_0_0_24;
   wire n_0_0_38;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_35;
   wire n_0_0_6;
   wire n_0_0_27;
   wire n_0_0_41;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_47;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_16;
   wire n_0_0_22;
   wire n_0_0_52;
   wire n_0_0_28;
   wire n_0_0_56;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_60;
   wire n_0_0_36;
   wire n_0_0_40;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_51;
   wire n_0_0_54;
   wire n_0_0_33;
   wire n_0_0_57;
   wire n_0_0_59;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_17;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_70;
   wire n_0_0_73;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_72;
   wire n_0_0_69;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_34;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_39;
   wire n_0_0_71;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;

   OAI22_X1 i_0_0_0 (.A1(A[0]), .A2(n_0_0_69), .B1(n_0_0_72), .B2(B[0]), 
      .ZN(result[0]));
   XOR2_X1 i_0_0_1 (.A(n_0_0_1), .B(n_0_0_0), .Z(result[1]));
   OAI221_X1 i_0_0_2 (.A(B[0]), .B1(n_0_0_72), .B2(n_0_0_71), .C1(A[0]), 
      .C2(is_subtract), .ZN(n_0_0_0));
   OAI22_X1 i_0_0_3 (.A1(n_0_0_73), .A2(n_0_0_70), .B1(A[1]), .B2(B[1]), 
      .ZN(n_0_0_1));
   XOR2_X1 i_0_0_4 (.A(n_0_0_27), .B(n_0_0_2), .Z(result[2]));
   AOI21_X1 i_0_0_5 (.A(n_0_0_33), .B1(A[2]), .B2(n_0_0_34), .ZN(n_0_0_2));
   XNOR2_X1 i_0_0_6 (.A(n_0_0_35), .B(n_0_0_26), .ZN(result[3]));
   XNOR2_X1 i_0_0_7 (.A(n_0_0_25), .B(n_0_0_3), .ZN(result[4]));
   NAND2_X1 i_0_0_8 (.A1(n_0_0_38), .A2(n_0_0_37), .ZN(n_0_0_3));
   XOR2_X1 i_0_0_9 (.A(n_0_0_24), .B(n_0_0_4), .Z(result[5]));
   OAI21_X1 i_0_0_10 (.A(n_0_0_41), .B1(A[5]), .B2(n_0_0_42), .ZN(n_0_0_4));
   XOR2_X1 i_0_0_11 (.A(n_0_0_43), .B(n_0_0_23), .Z(result[6]));
   XNOR2_X1 i_0_0_12 (.A(n_0_0_46), .B(n_0_0_21), .ZN(result[7]));
   XNOR2_X1 i_0_0_13 (.A(n_0_0_20), .B(n_0_0_19), .ZN(result[8]));
   XOR2_X1 i_0_0_14 (.A(n_0_0_18), .B(n_0_0_17), .Z(result[9]));
   XOR2_X1 i_0_0_15 (.A(n_0_0_15), .B(n_0_0_5), .Z(result[10]));
   OAI21_X1 i_0_0_16 (.A(n_0_0_52), .B1(A[10]), .B2(n_0_0_53), .ZN(n_0_0_5));
   XNOR2_X1 i_0_0_17 (.A(n_0_0_55), .B(n_0_0_14), .ZN(result[11]));
   XNOR2_X1 i_0_0_18 (.A(n_0_0_13), .B(n_0_0_12), .ZN(result[12]));
   NAND2_X1 i_0_0_19 (.A1(A[4]), .A2(n_0_0_39), .ZN(n_0_0_37));
   XNOR2_X1 i_0_0_20 (.A(n_0_0_71), .B(B[5]), .ZN(n_0_0_42));
   XNOR2_X1 i_0_0_21 (.A(A[7]), .B(n_0_0_47), .ZN(n_0_0_46));
   XNOR2_X1 i_0_0_22 (.A(is_subtract), .B(B[9]), .ZN(n_0_0_50));
   XNOR2_X1 i_0_0_23 (.A(n_0_0_71), .B(B[10]), .ZN(n_0_0_53));
   XNOR2_X1 i_0_0_24 (.A(A[11]), .B(n_0_0_56), .ZN(n_0_0_55));
   NAND2_X1 i_0_0_25 (.A1(A[13]), .A2(n_0_0_60), .ZN(n_0_0_58));
   XNOR2_X1 i_0_0_26 (.A(n_0_0_71), .B(B[14]), .ZN(n_0_0_63));
   XNOR2_X1 i_0_0_27 (.A(n_0_0_71), .B(B[15]), .ZN(n_0_0_68));
   AND2_X1 i_0_0_28 (.A1(n_0_0_54), .A2(n_0_0_82), .ZN(n_0_0_12));
   INV_X1 i_0_0_29 (.A(n_0_0_83), .ZN(n_0_0_13));
   NOR2_X1 i_0_0_30 (.A1(n_0_0_87), .A2(n_0_0_28), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_31 (.A1(n_0_0_89), .A2(n_0_0_88), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_32 (.A(n_0_0_94), .B1(n_0_0_20), .B2(n_0_0_132), .ZN(n_0_0_18));
   AND2_X1 i_0_0_33 (.A1(n_0_0_11), .A2(n_0_0_94), .ZN(n_0_0_19));
   INV_X1 i_0_0_34 (.A(n_0_0_95), .ZN(n_0_0_23));
   AND2_X1 i_0_0_35 (.A1(n_0_0_7), .A2(n_0_0_128), .ZN(n_0_0_43));
   INV_X1 i_0_0_36 (.A(n_0_0_96), .ZN(n_0_0_24));
   INV_X1 i_0_0_37 (.A(n_0_0_51), .ZN(n_0_0_38));
   INV_X1 i_0_0_38 (.A(n_0_0_49), .ZN(n_0_0_25));
   INV_X1 i_0_0_39 (.A(n_0_0_48), .ZN(n_0_0_26));
   NOR2_X1 i_0_0_40 (.A1(n_0_0_6), .A2(n_0_0_118), .ZN(n_0_0_35));
   INV_X1 i_0_0_41 (.A(n_0_0_45), .ZN(n_0_0_6));
   INV_X1 i_0_0_42 (.A(n_0_0_44), .ZN(n_0_0_27));
   NAND2_X1 i_0_0_43 (.A1(n_0_0_42), .A2(A[5]), .ZN(n_0_0_41));
   OR2_X1 i_0_0_44 (.A1(n_0_0_8), .A2(A[6]), .ZN(n_0_0_7));
   XNOR2_X1 i_0_0_45 (.A(n_0_0_71), .B(B[6]), .ZN(n_0_0_8));
   NAND2_X1 i_0_0_46 (.A1(n_0_0_47), .A2(A[7]), .ZN(n_0_0_9));
   INV_X1 i_0_0_47 (.A(n_0_0_10), .ZN(n_0_0_47));
   XNOR2_X1 i_0_0_48 (.A(is_subtract), .B(B[7]), .ZN(n_0_0_10));
   OR2_X1 i_0_0_49 (.A1(n_0_0_16), .A2(A[8]), .ZN(n_0_0_11));
   XNOR2_X1 i_0_0_50 (.A(n_0_0_71), .B(B[8]), .ZN(n_0_0_16));
   INV_X1 i_0_0_51 (.A(A[9]), .ZN(n_0_0_22));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_53), .A2(A[10]), .ZN(n_0_0_52));
   NOR2_X1 i_0_0_53 (.A1(n_0_0_53), .A2(A[10]), .ZN(n_0_0_28));
   INV_X1 i_0_0_54 (.A(n_0_0_29), .ZN(n_0_0_56));
   XNOR2_X1 i_0_0_55 (.A(is_subtract), .B(B[11]), .ZN(n_0_0_29));
   INV_X1 i_0_0_56 (.A(n_0_0_31), .ZN(n_0_0_30));
   XNOR2_X1 i_0_0_57 (.A(n_0_0_71), .B(B[12]), .ZN(n_0_0_31));
   INV_X1 i_0_0_58 (.A(A[12]), .ZN(n_0_0_32));
   INV_X1 i_0_0_59 (.A(n_0_0_36), .ZN(n_0_0_60));
   XNOR2_X1 i_0_0_60 (.A(is_subtract), .B(B[13]), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_61 (.A1(n_0_0_63), .A2(A[14]), .ZN(n_0_0_40));
   NAND2_X1 i_0_0_62 (.A1(n_0_0_100), .A2(n_0_0_107), .ZN(n_0_0_44));
   INV_X1 i_0_0_63 (.A(n_0_0_117), .ZN(n_0_0_45));
   NAND2_X1 i_0_0_64 (.A1(n_0_0_99), .A2(n_0_0_114), .ZN(n_0_0_48));
   NOR2_X1 i_0_0_65 (.A1(n_0_0_98), .A2(n_0_0_118), .ZN(n_0_0_49));
   INV_X1 i_0_0_66 (.A(n_0_0_122), .ZN(n_0_0_51));
   INV_X1 i_0_0_67 (.A(n_0_0_134), .ZN(n_0_0_54));
   INV_X1 i_0_0_68 (.A(n_0_0_112), .ZN(n_0_0_33));
   NAND2_X1 i_0_0_69 (.A1(n_0_0_78), .A2(n_0_0_140), .ZN(negative));
   NOR2_X1 i_0_0_70 (.A1(n_0_0_57), .A2(n_0_0_142), .ZN(carry));
   NOR2_X1 i_0_0_71 (.A1(n_0_0_61), .A2(n_0_0_57), .ZN(overflow_flag));
   AOI21_X1 i_0_0_72 (.A(n_0_0_59), .B1(n_0_0_80), .B2(n_0_0_137), .ZN(n_0_0_57));
   INV_X1 i_0_0_73 (.A(n_0_0_140), .ZN(n_0_0_59));
   INV_X1 i_0_0_74 (.A(n_0_0_62), .ZN(n_0_0_61));
   NAND3_X1 i_0_0_75 (.A1(n_0_0_80), .A2(n_0_0_141), .A3(n_0_0_137), .ZN(
      n_0_0_62));
   INV_X1 i_0_0_77 (.A(n_0_0_64), .ZN(result[13]));
   XNOR2_X1 i_0_0_82 (.A(n_0_0_81), .B(n_0_0_65), .ZN(n_0_0_64));
   OAI21_X1 i_0_0_86 (.A(n_0_0_58), .B1(n_0_0_60), .B2(A[13]), .ZN(n_0_0_65));
   INV_X1 i_0_0_76 (.A(n_0_0_66), .ZN(result[14]));
   NAND2_X1 i_0_0_78 (.A1(n_0_0_67), .A2(n_0_0_75), .ZN(n_0_0_66));
   NAND3_X1 i_0_0_79 (.A1(n_0_0_74), .A2(n_0_0_40), .A3(n_0_0_137), .ZN(n_0_0_67));
   OAI21_X1 i_0_0_80 (.A(n_0_0_136), .B1(n_0_0_81), .B2(n_0_0_135), .ZN(n_0_0_74));
   OAI211_X1 i_0_0_81 (.A(n_0_0_136), .B(n_0_0_76), .C1(n_0_0_81), .C2(n_0_0_135), 
      .ZN(n_0_0_75));
   NAND2_X1 i_0_0_83 (.A1(n_0_0_137), .A2(n_0_0_40), .ZN(n_0_0_76));
   NAND2_X1 i_0_0_84 (.A1(n_0_0_78), .A2(n_0_0_77), .ZN(result[15]));
   NAND3_X1 i_0_0_85 (.A1(n_0_0_80), .A2(n_0_0_139), .A3(n_0_0_137), .ZN(
      n_0_0_77));
   NAND2_X1 i_0_0_87 (.A1(n_0_0_79), .A2(n_0_0_138), .ZN(n_0_0_78));
   NAND2_X1 i_0_0_88 (.A1(n_0_0_80), .A2(n_0_0_137), .ZN(n_0_0_79));
   OAI211_X1 i_0_0_89 (.A(n_0_0_40), .B(n_0_0_136), .C1(n_0_0_81), .C2(n_0_0_135), 
      .ZN(n_0_0_80));
   AOI21_X1 i_0_0_90 (.A(n_0_0_134), .B1(n_0_0_83), .B2(n_0_0_82), .ZN(n_0_0_81));
   NAND2_X1 i_0_0_91 (.A1(n_0_0_30), .A2(n_0_0_32), .ZN(n_0_0_82));
   OAI21_X1 i_0_0_92 (.A(n_0_0_84), .B1(n_0_0_87), .B2(n_0_0_85), .ZN(n_0_0_83));
   NAND2_X1 i_0_0_93 (.A1(n_0_0_56), .A2(A[11]), .ZN(n_0_0_84));
   INV_X1 i_0_0_94 (.A(n_0_0_86), .ZN(n_0_0_85));
   NOR2_X1 i_0_0_95 (.A1(n_0_0_55), .A2(n_0_0_28), .ZN(n_0_0_86));
   AOI21_X1 i_0_0_96 (.A(n_0_0_133), .B1(n_0_0_89), .B2(n_0_0_88), .ZN(n_0_0_87));
   NAND2_X1 i_0_0_97 (.A1(n_0_0_50), .A2(n_0_0_22), .ZN(n_0_0_88));
   OAI21_X1 i_0_0_98 (.A(n_0_0_90), .B1(n_0_0_20), .B2(n_0_0_132), .ZN(n_0_0_89));
   INV_X1 i_0_0_99 (.A(n_0_0_91), .ZN(n_0_0_90));
   NAND2_X1 i_0_0_100 (.A1(n_0_0_17), .A2(n_0_0_94), .ZN(n_0_0_91));
   INV_X1 i_0_0_101 (.A(n_0_0_92), .ZN(n_0_0_17));
   XNOR2_X1 i_0_0_102 (.A(n_0_0_50), .B(n_0_0_93), .ZN(n_0_0_92));
   INV_X1 i_0_0_103 (.A(A[9]), .ZN(n_0_0_93));
   NAND2_X1 i_0_0_104 (.A1(n_0_0_16), .A2(A[8]), .ZN(n_0_0_94));
   AOI21_X1 i_0_0_105 (.A(n_0_0_130), .B1(n_0_0_131), .B2(n_0_0_21), .ZN(
      n_0_0_20));
   OAI21_X1 i_0_0_106 (.A(n_0_0_128), .B1(n_0_0_95), .B2(n_0_0_129), .ZN(
      n_0_0_21));
   AOI21_X1 i_0_0_107 (.A(n_0_0_127), .B1(n_0_0_96), .B2(n_0_0_126), .ZN(
      n_0_0_95));
   NAND2_X1 i_0_0_108 (.A1(n_0_0_97), .A2(n_0_0_125), .ZN(n_0_0_96));
   OAI21_X1 i_0_0_109 (.A(n_0_0_122), .B1(n_0_0_98), .B2(n_0_0_118), .ZN(
      n_0_0_97));
   AOI21_X1 i_0_0_110 (.A(n_0_0_117), .B1(n_0_0_99), .B2(n_0_0_114), .ZN(
      n_0_0_98));
   NAND3_X1 i_0_0_111 (.A1(n_0_0_107), .A2(n_0_0_100), .A3(n_0_0_112), .ZN(
      n_0_0_99));
   INV_X1 i_0_0_112 (.A(n_0_0_101), .ZN(n_0_0_100));
   NAND2_X1 i_0_0_113 (.A1(n_0_0_102), .A2(n_0_0_106), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_114 (.A1(n_0_0_105), .A2(n_0_0_103), .ZN(n_0_0_102));
   INV_X1 i_0_0_115 (.A(n_0_0_104), .ZN(n_0_0_103));
   NAND2_X1 i_0_0_116 (.A1(is_subtract), .A2(B[1]), .ZN(n_0_0_104));
   OAI21_X1 i_0_0_117 (.A(A[1]), .B1(n_0_0_69), .B2(A[0]), .ZN(n_0_0_105));
   NAND3_X1 i_0_0_118 (.A1(n_0_0_73), .A2(n_0_0_72), .A3(B[0]), .ZN(n_0_0_106));
   OAI21_X1 i_0_0_119 (.A(n_0_0_108), .B1(n_0_0_110), .B2(n_0_0_69), .ZN(
      n_0_0_107));
   INV_X1 i_0_0_120 (.A(n_0_0_109), .ZN(n_0_0_108));
   OAI21_X1 i_0_0_121 (.A(n_0_0_71), .B1(n_0_0_73), .B2(n_0_0_70), .ZN(n_0_0_109));
   INV_X1 i_0_0_122 (.A(B[1]), .ZN(n_0_0_70));
   INV_X1 i_0_0_123 (.A(A[1]), .ZN(n_0_0_73));
   AOI21_X1 i_0_0_124 (.A(B[1]), .B1(n_0_0_111), .B2(A[1]), .ZN(n_0_0_110));
   NAND2_X1 i_0_0_125 (.A1(n_0_0_72), .A2(B[0]), .ZN(n_0_0_111));
   INV_X1 i_0_0_126 (.A(A[0]), .ZN(n_0_0_72));
   INV_X1 i_0_0_127 (.A(B[0]), .ZN(n_0_0_69));
   NAND3_X1 i_0_0_128 (.A1(n_0_0_116), .A2(n_0_0_115), .A3(n_0_0_113), .ZN(
      n_0_0_112));
   INV_X1 i_0_0_129 (.A(A[2]), .ZN(n_0_0_113));
   NAND2_X1 i_0_0_130 (.A1(n_0_0_34), .A2(A[2]), .ZN(n_0_0_114));
   NAND2_X1 i_0_0_131 (.A1(n_0_0_116), .A2(n_0_0_115), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_132 (.A1(n_0_0_71), .A2(B[2]), .ZN(n_0_0_115));
   OR2_X1 i_0_0_133 (.A1(n_0_0_71), .A2(B[2]), .ZN(n_0_0_116));
   NOR2_X1 i_0_0_134 (.A1(n_0_0_120), .A2(A[3]), .ZN(n_0_0_117));
   INV_X1 i_0_0_135 (.A(n_0_0_119), .ZN(n_0_0_118));
   NAND2_X1 i_0_0_136 (.A1(n_0_0_120), .A2(A[3]), .ZN(n_0_0_119));
   INV_X1 i_0_0_137 (.A(n_0_0_121), .ZN(n_0_0_120));
   XNOR2_X1 i_0_0_138 (.A(is_subtract), .B(B[3]), .ZN(n_0_0_121));
   NAND2_X1 i_0_0_139 (.A1(n_0_0_123), .A2(n_0_0_124), .ZN(n_0_0_122));
   INV_X1 i_0_0_140 (.A(n_0_0_39), .ZN(n_0_0_123));
   INV_X1 i_0_0_141 (.A(A[4]), .ZN(n_0_0_124));
   NAND2_X1 i_0_0_142 (.A1(n_0_0_39), .A2(A[4]), .ZN(n_0_0_125));
   XNOR2_X1 i_0_0_143 (.A(n_0_0_71), .B(B[4]), .ZN(n_0_0_39));
   INV_X1 i_0_0_144 (.A(is_subtract), .ZN(n_0_0_71));
   OR2_X1 i_0_0_145 (.A1(n_0_0_42), .A2(A[5]), .ZN(n_0_0_126));
   INV_X1 i_0_0_146 (.A(n_0_0_41), .ZN(n_0_0_127));
   NAND2_X1 i_0_0_147 (.A1(n_0_0_8), .A2(A[6]), .ZN(n_0_0_128));
   INV_X1 i_0_0_148 (.A(n_0_0_7), .ZN(n_0_0_129));
   INV_X1 i_0_0_149 (.A(n_0_0_9), .ZN(n_0_0_130));
   INV_X1 i_0_0_150 (.A(n_0_0_46), .ZN(n_0_0_131));
   INV_X1 i_0_0_151 (.A(n_0_0_11), .ZN(n_0_0_132));
   INV_X1 i_0_0_152 (.A(n_0_0_52), .ZN(n_0_0_133));
   NOR2_X1 i_0_0_153 (.A1(n_0_0_30), .A2(n_0_0_32), .ZN(n_0_0_134));
   NOR2_X1 i_0_0_154 (.A1(n_0_0_60), .A2(A[13]), .ZN(n_0_0_135));
   NAND2_X1 i_0_0_155 (.A1(n_0_0_60), .A2(A[13]), .ZN(n_0_0_136));
   OR2_X1 i_0_0_156 (.A1(n_0_0_63), .A2(A[14]), .ZN(n_0_0_137));
   INV_X1 i_0_0_157 (.A(n_0_0_139), .ZN(n_0_0_138));
   NAND2_X1 i_0_0_158 (.A1(n_0_0_141), .A2(n_0_0_140), .ZN(n_0_0_139));
   NAND2_X1 i_0_0_159 (.A1(n_0_0_68), .A2(A[15]), .ZN(n_0_0_140));
   INV_X1 i_0_0_160 (.A(n_0_0_142), .ZN(n_0_0_141));
   NOR2_X1 i_0_0_161 (.A1(n_0_0_68), .A2(A[15]), .ZN(n_0_0_142));
endmodule
