/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 20:07:21 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3911429606 */

module memory_manager(clk, reset, store1, store2, write, temp1, temp2, data1, 
      data2, select);
   input clk;
   input reset;
   input store1;
   input store2;
   output write;
   output [31:0]temp1;
   output [31:0]temp2;
   input [31:0]data1;
   input [31:0]data2;
   output [1:0]select;

   wire counter;
   wire wait2;
   wire wait1;
   wire n_0_2;
   wire n_0_0;
   wire n_0_0_0;
   wire n_0_1;
   wire n_0_0_1;
   wire n_0_4;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_5;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_6;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_7;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_9;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_10;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_71;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_70;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_69;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_68;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_67;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_66;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_65;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_64;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_63;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_62;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_61;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_60;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_59;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_58;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_57;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_56;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_55;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_53;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_52;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_51;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_50;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_49;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_48;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_47;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_46;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_45;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_44;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_43;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_42;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_41;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_40;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_39;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_38;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_37;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_36;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_35;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_34;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_33;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_32;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_31;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_30;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_29;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_28;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_27;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_26;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_25;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_24;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_23;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_22;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_21;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_20;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_19;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_18;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_17;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_16;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_15;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_14;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_11;
   wire n_0_0_143;
   wire n_0_12;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_8;
   wire n_0_13;
   wire n_0_3;
   wire n_0_0_7;
   wire n_0_0_8;

   DFFR_X1 counter_reg (.D(n_0_13), .RN(n_0_8), .CK(clk), .Q(counter), .QN());
   DFF_X1 \select_reg[1]  (.D(n_0_12), .CK(n_0_2), .Q(select[1]), .QN());
   DFF_X1 \select_reg[0]  (.D(n_0_11), .CK(n_0_2), .Q(select[0]), .QN());
   DFF_X1 \temp2_reg[31]  (.D(n_0_14), .CK(n_0_2), .Q(temp2[31]), .QN());
   DFF_X1 \temp2_reg[30]  (.D(n_0_15), .CK(n_0_2), .Q(temp2[30]), .QN());
   DFF_X1 \temp2_reg[29]  (.D(n_0_16), .CK(n_0_2), .Q(temp2[29]), .QN());
   DFF_X1 \temp2_reg[28]  (.D(n_0_17), .CK(n_0_2), .Q(temp2[28]), .QN());
   DFF_X1 \temp2_reg[27]  (.D(n_0_18), .CK(n_0_2), .Q(temp2[27]), .QN());
   DFF_X1 \temp2_reg[26]  (.D(n_0_19), .CK(n_0_2), .Q(temp2[26]), .QN());
   DFF_X1 \temp2_reg[25]  (.D(n_0_20), .CK(n_0_2), .Q(temp2[25]), .QN());
   DFF_X1 \temp2_reg[24]  (.D(n_0_21), .CK(n_0_2), .Q(temp2[24]), .QN());
   DFF_X1 \temp2_reg[23]  (.D(n_0_22), .CK(n_0_2), .Q(temp2[23]), .QN());
   DFF_X1 \temp2_reg[22]  (.D(n_0_23), .CK(n_0_2), .Q(temp2[22]), .QN());
   DFF_X1 \temp2_reg[21]  (.D(n_0_24), .CK(n_0_2), .Q(temp2[21]), .QN());
   DFF_X1 \temp2_reg[20]  (.D(n_0_25), .CK(n_0_2), .Q(temp2[20]), .QN());
   DFF_X1 \temp2_reg[19]  (.D(n_0_26), .CK(n_0_2), .Q(temp2[19]), .QN());
   DFF_X1 \temp2_reg[18]  (.D(n_0_27), .CK(n_0_2), .Q(temp2[18]), .QN());
   DFF_X1 \temp2_reg[17]  (.D(n_0_28), .CK(n_0_2), .Q(temp2[17]), .QN());
   DFF_X1 \temp2_reg[16]  (.D(n_0_29), .CK(n_0_2), .Q(temp2[16]), .QN());
   DFF_X1 \temp2_reg[15]  (.D(n_0_30), .CK(n_0_2), .Q(temp2[15]), .QN());
   DFF_X1 \temp2_reg[14]  (.D(n_0_31), .CK(n_0_2), .Q(temp2[14]), .QN());
   DFF_X1 \temp2_reg[13]  (.D(n_0_32), .CK(n_0_2), .Q(temp2[13]), .QN());
   DFF_X1 \temp2_reg[12]  (.D(n_0_33), .CK(n_0_2), .Q(temp2[12]), .QN());
   DFF_X1 \temp2_reg[11]  (.D(n_0_34), .CK(n_0_2), .Q(temp2[11]), .QN());
   DFF_X1 \temp2_reg[10]  (.D(n_0_35), .CK(n_0_2), .Q(temp2[10]), .QN());
   DFF_X1 \temp2_reg[9]  (.D(n_0_36), .CK(n_0_2), .Q(temp2[9]), .QN());
   DFF_X1 \temp2_reg[8]  (.D(n_0_37), .CK(n_0_2), .Q(temp2[8]), .QN());
   DFF_X1 \temp2_reg[7]  (.D(n_0_38), .CK(n_0_2), .Q(temp2[7]), .QN());
   DFF_X1 \temp2_reg[6]  (.D(n_0_39), .CK(n_0_2), .Q(temp2[6]), .QN());
   DFF_X1 \temp2_reg[5]  (.D(n_0_40), .CK(n_0_2), .Q(temp2[5]), .QN());
   DFF_X1 \temp2_reg[4]  (.D(n_0_41), .CK(n_0_2), .Q(temp2[4]), .QN());
   DFF_X1 \temp2_reg[3]  (.D(n_0_42), .CK(n_0_2), .Q(temp2[3]), .QN());
   DFF_X1 \temp2_reg[2]  (.D(n_0_43), .CK(n_0_2), .Q(temp2[2]), .QN());
   DFF_X1 \temp2_reg[1]  (.D(n_0_44), .CK(n_0_2), .Q(temp2[1]), .QN());
   DFF_X1 \temp2_reg[0]  (.D(n_0_45), .CK(n_0_2), .Q(temp2[0]), .QN());
   DFF_X1 \temp1_reg[31]  (.D(n_0_46), .CK(n_0_2), .Q(temp1[31]), .QN());
   DFF_X1 \temp1_reg[30]  (.D(n_0_47), .CK(n_0_2), .Q(temp1[30]), .QN());
   DFF_X1 \temp1_reg[29]  (.D(n_0_48), .CK(n_0_2), .Q(temp1[29]), .QN());
   DFF_X1 \temp1_reg[28]  (.D(n_0_49), .CK(n_0_2), .Q(temp1[28]), .QN());
   DFF_X1 \temp1_reg[27]  (.D(n_0_50), .CK(n_0_2), .Q(temp1[27]), .QN());
   DFF_X1 \temp1_reg[26]  (.D(n_0_51), .CK(n_0_2), .Q(temp1[26]), .QN());
   DFF_X1 \temp1_reg[25]  (.D(n_0_52), .CK(n_0_2), .Q(temp1[25]), .QN());
   DFF_X1 \temp1_reg[24]  (.D(n_0_53), .CK(n_0_2), .Q(temp1[24]), .QN());
   DFF_X1 \temp1_reg[23]  (.D(n_0_54), .CK(n_0_2), .Q(temp1[23]), .QN());
   DFF_X1 \temp1_reg[22]  (.D(n_0_55), .CK(n_0_2), .Q(temp1[22]), .QN());
   DFF_X1 \temp1_reg[21]  (.D(n_0_56), .CK(n_0_2), .Q(temp1[21]), .QN());
   DFF_X1 \temp1_reg[20]  (.D(n_0_57), .CK(n_0_2), .Q(temp1[20]), .QN());
   DFF_X1 \temp1_reg[19]  (.D(n_0_58), .CK(n_0_2), .Q(temp1[19]), .QN());
   DFF_X1 \temp1_reg[18]  (.D(n_0_59), .CK(n_0_2), .Q(temp1[18]), .QN());
   DFF_X1 \temp1_reg[17]  (.D(n_0_60), .CK(n_0_2), .Q(temp1[17]), .QN());
   DFF_X1 \temp1_reg[16]  (.D(n_0_61), .CK(n_0_2), .Q(temp1[16]), .QN());
   DFF_X1 \temp1_reg[15]  (.D(n_0_62), .CK(n_0_2), .Q(temp1[15]), .QN());
   DFF_X1 \temp1_reg[14]  (.D(n_0_63), .CK(n_0_2), .Q(temp1[14]), .QN());
   DFF_X1 \temp1_reg[13]  (.D(n_0_64), .CK(n_0_2), .Q(temp1[13]), .QN());
   DFF_X1 \temp1_reg[12]  (.D(n_0_65), .CK(n_0_2), .Q(temp1[12]), .QN());
   DFF_X1 \temp1_reg[11]  (.D(n_0_66), .CK(n_0_2), .Q(temp1[11]), .QN());
   DFF_X1 \temp1_reg[10]  (.D(n_0_67), .CK(n_0_2), .Q(temp1[10]), .QN());
   DFF_X1 \temp1_reg[9]  (.D(n_0_68), .CK(n_0_2), .Q(temp1[9]), .QN());
   DFF_X1 \temp1_reg[8]  (.D(n_0_69), .CK(n_0_2), .Q(temp1[8]), .QN());
   DFF_X1 \temp1_reg[7]  (.D(n_0_70), .CK(n_0_2), .Q(temp1[7]), .QN());
   DFF_X1 \temp1_reg[6]  (.D(n_0_71), .CK(n_0_2), .Q(temp1[6]), .QN());
   DFF_X1 \temp1_reg[5]  (.D(n_0_10), .CK(n_0_2), .Q(temp1[5]), .QN());
   DFF_X1 \temp1_reg[4]  (.D(n_0_9), .CK(n_0_2), .Q(temp1[4]), .QN());
   DFF_X1 \temp1_reg[3]  (.D(n_0_7), .CK(n_0_2), .Q(temp1[3]), .QN());
   DFF_X1 \temp1_reg[2]  (.D(n_0_6), .CK(n_0_2), .Q(temp1[2]), .QN());
   DFF_X1 \temp1_reg[1]  (.D(n_0_5), .CK(n_0_2), .Q(temp1[1]), .QN());
   DFF_X1 \temp1_reg[0]  (.D(n_0_4), .CK(n_0_2), .Q(temp1[0]), .QN());
   DFF_X1 write_reg (.D(n_0_3), .CK(n_0_2), .Q(write), .QN());
   DFF_X1 wait2_reg (.D(n_0_1), .CK(n_0_2), .Q(wait2), .QN());
   DFF_X1 wait1_reg (.D(n_0_0), .CK(n_0_2), .Q(wait1), .QN());
   INV_X1 i_0_0_84 (.A(clk), .ZN(n_0_2));
   NAND2_X1 i_0_0_0 (.A1(n_0_0_75), .A2(n_0_0_0), .ZN(n_0_0));
   NAND3_X1 i_0_0_1 (.A1(n_0_8), .A2(counter), .A3(wait1), .ZN(n_0_0_0));
   NAND2_X1 i_0_0_2 (.A1(n_0_0_139), .A2(n_0_0_1), .ZN(n_0_1));
   NAND3_X1 i_0_0_3 (.A1(n_0_8), .A2(n_0_13), .A3(wait2), .ZN(n_0_0_1));
   NAND2_X1 i_0_0_12 (.A1(n_0_0_9), .A2(n_0_0_10), .ZN(n_0_4));
   NAND3_X1 i_0_0_13 (.A1(n_0_0_72), .A2(data1[0]), .A3(store1), .ZN(n_0_0_9));
   NAND2_X1 i_0_0_14 (.A1(n_0_0_75), .A2(temp1[0]), .ZN(n_0_0_10));
   NAND2_X1 i_0_0_15 (.A1(n_0_0_11), .A2(n_0_0_12), .ZN(n_0_5));
   NAND3_X1 i_0_0_16 (.A1(n_0_0_72), .A2(data1[1]), .A3(store1), .ZN(n_0_0_11));
   NAND2_X1 i_0_0_17 (.A1(n_0_0_75), .A2(temp1[1]), .ZN(n_0_0_12));
   NAND2_X1 i_0_0_18 (.A1(n_0_0_13), .A2(n_0_0_14), .ZN(n_0_6));
   NAND3_X1 i_0_0_19 (.A1(n_0_0_72), .A2(data1[2]), .A3(store1), .ZN(n_0_0_13));
   NAND2_X1 i_0_0_20 (.A1(n_0_0_75), .A2(temp1[2]), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_21 (.A1(n_0_0_15), .A2(n_0_0_16), .ZN(n_0_7));
   NAND3_X1 i_0_0_22 (.A1(n_0_0_72), .A2(data1[3]), .A3(store1), .ZN(n_0_0_15));
   NAND2_X1 i_0_0_23 (.A1(n_0_0_75), .A2(temp1[3]), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_24 (.A1(n_0_0_17), .A2(n_0_0_18), .ZN(n_0_9));
   NAND3_X1 i_0_0_25 (.A1(n_0_0_72), .A2(data1[4]), .A3(store1), .ZN(n_0_0_17));
   NAND2_X1 i_0_0_26 (.A1(n_0_0_75), .A2(temp1[4]), .ZN(n_0_0_18));
   NAND2_X1 i_0_0_27 (.A1(n_0_0_19), .A2(n_0_0_20), .ZN(n_0_10));
   NAND3_X1 i_0_0_28 (.A1(n_0_0_72), .A2(data1[5]), .A3(store1), .ZN(n_0_0_19));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_75), .A2(temp1[5]), .ZN(n_0_0_20));
   NAND2_X1 i_0_0_30 (.A1(n_0_0_21), .A2(n_0_0_22), .ZN(n_0_71));
   NAND3_X1 i_0_0_31 (.A1(n_0_0_72), .A2(data1[6]), .A3(store1), .ZN(n_0_0_21));
   NAND2_X1 i_0_0_32 (.A1(n_0_0_75), .A2(temp1[6]), .ZN(n_0_0_22));
   NAND2_X1 i_0_0_33 (.A1(n_0_0_23), .A2(n_0_0_24), .ZN(n_0_70));
   NAND3_X1 i_0_0_34 (.A1(n_0_0_72), .A2(data1[7]), .A3(store1), .ZN(n_0_0_23));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_75), .A2(temp1[7]), .ZN(n_0_0_24));
   NAND2_X1 i_0_0_36 (.A1(n_0_0_25), .A2(n_0_0_26), .ZN(n_0_69));
   NAND3_X1 i_0_0_37 (.A1(n_0_0_72), .A2(data1[8]), .A3(store1), .ZN(n_0_0_25));
   NAND2_X1 i_0_0_38 (.A1(n_0_0_75), .A2(temp1[8]), .ZN(n_0_0_26));
   NAND2_X1 i_0_0_39 (.A1(n_0_0_27), .A2(n_0_0_28), .ZN(n_0_68));
   NAND3_X1 i_0_0_40 (.A1(n_0_0_72), .A2(data1[9]), .A3(store1), .ZN(n_0_0_27));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_75), .A2(temp1[9]), .ZN(n_0_0_28));
   NAND2_X1 i_0_0_42 (.A1(n_0_0_29), .A2(n_0_0_30), .ZN(n_0_67));
   NAND3_X1 i_0_0_43 (.A1(n_0_0_72), .A2(data1[10]), .A3(store1), .ZN(n_0_0_29));
   NAND2_X1 i_0_0_44 (.A1(n_0_0_75), .A2(temp1[10]), .ZN(n_0_0_30));
   NAND2_X1 i_0_0_45 (.A1(n_0_0_31), .A2(n_0_0_32), .ZN(n_0_66));
   NAND3_X1 i_0_0_46 (.A1(n_0_0_72), .A2(data1[11]), .A3(store1), .ZN(n_0_0_31));
   NAND2_X1 i_0_0_47 (.A1(n_0_0_75), .A2(temp1[11]), .ZN(n_0_0_32));
   NAND2_X1 i_0_0_48 (.A1(n_0_0_33), .A2(n_0_0_34), .ZN(n_0_65));
   NAND3_X1 i_0_0_49 (.A1(n_0_0_72), .A2(data1[12]), .A3(store1), .ZN(n_0_0_33));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_75), .A2(temp1[12]), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_51 (.A1(n_0_0_35), .A2(n_0_0_36), .ZN(n_0_64));
   NAND3_X1 i_0_0_52 (.A1(n_0_0_72), .A2(data1[13]), .A3(store1), .ZN(n_0_0_35));
   NAND2_X1 i_0_0_53 (.A1(n_0_0_75), .A2(temp1[13]), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_54 (.A1(n_0_0_37), .A2(n_0_0_38), .ZN(n_0_63));
   NAND3_X1 i_0_0_55 (.A1(n_0_0_72), .A2(data1[14]), .A3(store1), .ZN(n_0_0_37));
   NAND2_X1 i_0_0_56 (.A1(n_0_0_75), .A2(temp1[14]), .ZN(n_0_0_38));
   NAND2_X1 i_0_0_57 (.A1(n_0_0_39), .A2(n_0_0_40), .ZN(n_0_62));
   NAND3_X1 i_0_0_58 (.A1(n_0_0_72), .A2(data1[15]), .A3(store1), .ZN(n_0_0_39));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_75), .A2(temp1[15]), .ZN(n_0_0_40));
   NAND2_X1 i_0_0_60 (.A1(n_0_0_41), .A2(n_0_0_42), .ZN(n_0_61));
   NAND3_X1 i_0_0_61 (.A1(n_0_0_72), .A2(data1[16]), .A3(store1), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_62 (.A1(n_0_0_75), .A2(temp1[16]), .ZN(n_0_0_42));
   NAND2_X1 i_0_0_63 (.A1(n_0_0_43), .A2(n_0_0_44), .ZN(n_0_60));
   NAND3_X1 i_0_0_64 (.A1(n_0_0_72), .A2(data1[17]), .A3(store1), .ZN(n_0_0_43));
   NAND2_X1 i_0_0_65 (.A1(n_0_0_75), .A2(temp1[17]), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_66 (.A1(n_0_0_45), .A2(n_0_0_46), .ZN(n_0_59));
   NAND3_X1 i_0_0_67 (.A1(n_0_0_72), .A2(data1[18]), .A3(store1), .ZN(n_0_0_45));
   NAND2_X1 i_0_0_68 (.A1(n_0_0_75), .A2(temp1[18]), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_69 (.A1(n_0_0_47), .A2(n_0_0_48), .ZN(n_0_58));
   NAND3_X1 i_0_0_70 (.A1(n_0_0_72), .A2(data1[19]), .A3(store1), .ZN(n_0_0_47));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_75), .A2(temp1[19]), .ZN(n_0_0_48));
   NAND2_X1 i_0_0_72 (.A1(n_0_0_49), .A2(n_0_0_50), .ZN(n_0_57));
   NAND3_X1 i_0_0_73 (.A1(n_0_0_72), .A2(data1[20]), .A3(store1), .ZN(n_0_0_49));
   NAND2_X1 i_0_0_74 (.A1(n_0_0_75), .A2(temp1[20]), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_75 (.A1(n_0_0_51), .A2(n_0_0_52), .ZN(n_0_56));
   NAND3_X1 i_0_0_76 (.A1(n_0_0_72), .A2(data1[21]), .A3(store1), .ZN(n_0_0_51));
   NAND2_X1 i_0_0_77 (.A1(n_0_0_75), .A2(temp1[21]), .ZN(n_0_0_52));
   NAND2_X1 i_0_0_78 (.A1(n_0_0_53), .A2(n_0_0_54), .ZN(n_0_55));
   NAND3_X1 i_0_0_79 (.A1(n_0_0_72), .A2(data1[22]), .A3(store1), .ZN(n_0_0_53));
   NAND2_X1 i_0_0_80 (.A1(n_0_0_75), .A2(temp1[22]), .ZN(n_0_0_54));
   NAND2_X1 i_0_0_81 (.A1(n_0_0_55), .A2(n_0_0_56), .ZN(n_0_54));
   NAND3_X1 i_0_0_82 (.A1(n_0_0_72), .A2(data1[23]), .A3(store1), .ZN(n_0_0_55));
   NAND2_X1 i_0_0_83 (.A1(n_0_0_75), .A2(temp1[23]), .ZN(n_0_0_56));
   NAND2_X1 i_0_0_85 (.A1(n_0_0_57), .A2(n_0_0_58), .ZN(n_0_53));
   NAND3_X1 i_0_0_86 (.A1(n_0_0_72), .A2(data1[24]), .A3(store1), .ZN(n_0_0_57));
   NAND2_X1 i_0_0_87 (.A1(n_0_0_75), .A2(temp1[24]), .ZN(n_0_0_58));
   NAND2_X1 i_0_0_88 (.A1(n_0_0_59), .A2(n_0_0_60), .ZN(n_0_52));
   NAND3_X1 i_0_0_89 (.A1(n_0_0_72), .A2(data1[25]), .A3(store1), .ZN(n_0_0_59));
   NAND2_X1 i_0_0_90 (.A1(n_0_0_75), .A2(temp1[25]), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_91 (.A1(n_0_0_61), .A2(n_0_0_62), .ZN(n_0_51));
   NAND3_X1 i_0_0_92 (.A1(n_0_0_72), .A2(data1[26]), .A3(store1), .ZN(n_0_0_61));
   NAND2_X1 i_0_0_93 (.A1(n_0_0_75), .A2(temp1[26]), .ZN(n_0_0_62));
   NAND2_X1 i_0_0_94 (.A1(n_0_0_63), .A2(n_0_0_64), .ZN(n_0_50));
   NAND3_X1 i_0_0_95 (.A1(n_0_0_72), .A2(data1[27]), .A3(store1), .ZN(n_0_0_63));
   NAND2_X1 i_0_0_96 (.A1(n_0_0_75), .A2(temp1[27]), .ZN(n_0_0_64));
   NAND2_X1 i_0_0_97 (.A1(n_0_0_65), .A2(n_0_0_66), .ZN(n_0_49));
   NAND3_X1 i_0_0_98 (.A1(n_0_0_72), .A2(data1[28]), .A3(store1), .ZN(n_0_0_65));
   NAND2_X1 i_0_0_99 (.A1(n_0_0_75), .A2(temp1[28]), .ZN(n_0_0_66));
   NAND2_X1 i_0_0_100 (.A1(n_0_0_67), .A2(n_0_0_68), .ZN(n_0_48));
   NAND3_X1 i_0_0_101 (.A1(n_0_0_72), .A2(data1[29]), .A3(store1), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_102 (.A1(n_0_0_75), .A2(temp1[29]), .ZN(n_0_0_68));
   NAND2_X1 i_0_0_103 (.A1(n_0_0_69), .A2(n_0_0_70), .ZN(n_0_47));
   NAND3_X1 i_0_0_104 (.A1(n_0_0_72), .A2(data1[30]), .A3(store1), .ZN(n_0_0_69));
   NAND2_X1 i_0_0_105 (.A1(n_0_0_75), .A2(temp1[30]), .ZN(n_0_0_70));
   NAND2_X1 i_0_0_106 (.A1(n_0_0_71), .A2(n_0_0_74), .ZN(n_0_46));
   NAND3_X1 i_0_0_107 (.A1(n_0_0_72), .A2(data1[31]), .A3(store1), .ZN(n_0_0_71));
   INV_X1 i_0_0_108 (.A(n_0_0_73), .ZN(n_0_0_72));
   OAI21_X1 i_0_0_109 (.A(n_0_8), .B1(counter), .B2(wait1), .ZN(n_0_0_73));
   NAND2_X1 i_0_0_110 (.A1(n_0_0_75), .A2(temp1[31]), .ZN(n_0_0_74));
   OAI211_X1 i_0_0_111 (.A(n_0_8), .B(store1), .C1(counter), .C2(wait1), 
      .ZN(n_0_0_75));
   OAI21_X1 i_0_0_112 (.A(n_0_0_76), .B1(n_0_0_77), .B2(n_0_0_139), .ZN(n_0_45));
   NAND2_X1 i_0_0_113 (.A1(n_0_0_139), .A2(temp2[0]), .ZN(n_0_0_76));
   INV_X1 i_0_0_114 (.A(data2[0]), .ZN(n_0_0_77));
   OAI21_X1 i_0_0_115 (.A(n_0_0_78), .B1(n_0_0_79), .B2(n_0_0_139), .ZN(n_0_44));
   NAND2_X1 i_0_0_116 (.A1(n_0_0_139), .A2(temp2[1]), .ZN(n_0_0_78));
   INV_X1 i_0_0_117 (.A(data2[1]), .ZN(n_0_0_79));
   OAI21_X1 i_0_0_118 (.A(n_0_0_80), .B1(n_0_0_81), .B2(n_0_0_139), .ZN(n_0_43));
   NAND2_X1 i_0_0_119 (.A1(n_0_0_139), .A2(temp2[2]), .ZN(n_0_0_80));
   INV_X1 i_0_0_120 (.A(data2[2]), .ZN(n_0_0_81));
   OAI21_X1 i_0_0_121 (.A(n_0_0_82), .B1(n_0_0_83), .B2(n_0_0_139), .ZN(n_0_42));
   NAND2_X1 i_0_0_122 (.A1(n_0_0_139), .A2(temp2[3]), .ZN(n_0_0_82));
   INV_X1 i_0_0_123 (.A(data2[3]), .ZN(n_0_0_83));
   OAI21_X1 i_0_0_124 (.A(n_0_0_84), .B1(n_0_0_85), .B2(n_0_0_139), .ZN(n_0_41));
   NAND2_X1 i_0_0_125 (.A1(n_0_0_139), .A2(temp2[4]), .ZN(n_0_0_84));
   INV_X1 i_0_0_126 (.A(data2[4]), .ZN(n_0_0_85));
   OAI21_X1 i_0_0_127 (.A(n_0_0_86), .B1(n_0_0_87), .B2(n_0_0_139), .ZN(n_0_40));
   NAND2_X1 i_0_0_128 (.A1(n_0_0_139), .A2(temp2[5]), .ZN(n_0_0_86));
   INV_X1 i_0_0_129 (.A(data2[5]), .ZN(n_0_0_87));
   OAI21_X1 i_0_0_130 (.A(n_0_0_88), .B1(n_0_0_89), .B2(n_0_0_139), .ZN(n_0_39));
   NAND2_X1 i_0_0_131 (.A1(n_0_0_139), .A2(temp2[6]), .ZN(n_0_0_88));
   INV_X1 i_0_0_132 (.A(data2[6]), .ZN(n_0_0_89));
   OAI21_X1 i_0_0_133 (.A(n_0_0_90), .B1(n_0_0_91), .B2(n_0_0_139), .ZN(n_0_38));
   NAND2_X1 i_0_0_134 (.A1(n_0_0_139), .A2(temp2[7]), .ZN(n_0_0_90));
   INV_X1 i_0_0_135 (.A(data2[7]), .ZN(n_0_0_91));
   OAI21_X1 i_0_0_136 (.A(n_0_0_92), .B1(n_0_0_93), .B2(n_0_0_139), .ZN(n_0_37));
   NAND2_X1 i_0_0_137 (.A1(n_0_0_139), .A2(temp2[8]), .ZN(n_0_0_92));
   INV_X1 i_0_0_138 (.A(data2[8]), .ZN(n_0_0_93));
   OAI21_X1 i_0_0_139 (.A(n_0_0_94), .B1(n_0_0_95), .B2(n_0_0_139), .ZN(n_0_36));
   NAND2_X1 i_0_0_140 (.A1(n_0_0_139), .A2(temp2[9]), .ZN(n_0_0_94));
   INV_X1 i_0_0_141 (.A(data2[9]), .ZN(n_0_0_95));
   OAI21_X1 i_0_0_142 (.A(n_0_0_96), .B1(n_0_0_97), .B2(n_0_0_139), .ZN(n_0_35));
   NAND2_X1 i_0_0_143 (.A1(n_0_0_139), .A2(temp2[10]), .ZN(n_0_0_96));
   INV_X1 i_0_0_144 (.A(data2[10]), .ZN(n_0_0_97));
   OAI21_X1 i_0_0_145 (.A(n_0_0_98), .B1(n_0_0_99), .B2(n_0_0_139), .ZN(n_0_34));
   NAND2_X1 i_0_0_146 (.A1(n_0_0_139), .A2(temp2[11]), .ZN(n_0_0_98));
   INV_X1 i_0_0_147 (.A(data2[11]), .ZN(n_0_0_99));
   OAI21_X1 i_0_0_148 (.A(n_0_0_100), .B1(n_0_0_101), .B2(n_0_0_139), .ZN(n_0_33));
   NAND2_X1 i_0_0_149 (.A1(n_0_0_139), .A2(temp2[12]), .ZN(n_0_0_100));
   INV_X1 i_0_0_150 (.A(data2[12]), .ZN(n_0_0_101));
   OAI21_X1 i_0_0_151 (.A(n_0_0_102), .B1(n_0_0_103), .B2(n_0_0_139), .ZN(n_0_32));
   NAND2_X1 i_0_0_152 (.A1(n_0_0_139), .A2(temp2[13]), .ZN(n_0_0_102));
   INV_X1 i_0_0_153 (.A(data2[13]), .ZN(n_0_0_103));
   OAI21_X1 i_0_0_154 (.A(n_0_0_104), .B1(n_0_0_105), .B2(n_0_0_139), .ZN(n_0_31));
   NAND2_X1 i_0_0_155 (.A1(n_0_0_139), .A2(temp2[14]), .ZN(n_0_0_104));
   INV_X1 i_0_0_156 (.A(data2[14]), .ZN(n_0_0_105));
   OAI21_X1 i_0_0_157 (.A(n_0_0_106), .B1(n_0_0_107), .B2(n_0_0_139), .ZN(n_0_30));
   NAND2_X1 i_0_0_158 (.A1(n_0_0_139), .A2(temp2[15]), .ZN(n_0_0_106));
   INV_X1 i_0_0_159 (.A(data2[15]), .ZN(n_0_0_107));
   OAI21_X1 i_0_0_160 (.A(n_0_0_108), .B1(n_0_0_109), .B2(n_0_0_139), .ZN(n_0_29));
   NAND2_X1 i_0_0_161 (.A1(n_0_0_139), .A2(temp2[16]), .ZN(n_0_0_108));
   INV_X1 i_0_0_162 (.A(data2[16]), .ZN(n_0_0_109));
   OAI21_X1 i_0_0_163 (.A(n_0_0_110), .B1(n_0_0_111), .B2(n_0_0_139), .ZN(n_0_28));
   NAND2_X1 i_0_0_164 (.A1(n_0_0_139), .A2(temp2[17]), .ZN(n_0_0_110));
   INV_X1 i_0_0_165 (.A(data2[17]), .ZN(n_0_0_111));
   OAI21_X1 i_0_0_166 (.A(n_0_0_112), .B1(n_0_0_113), .B2(n_0_0_139), .ZN(n_0_27));
   NAND2_X1 i_0_0_167 (.A1(n_0_0_139), .A2(temp2[18]), .ZN(n_0_0_112));
   INV_X1 i_0_0_168 (.A(data2[18]), .ZN(n_0_0_113));
   OAI21_X1 i_0_0_169 (.A(n_0_0_114), .B1(n_0_0_115), .B2(n_0_0_139), .ZN(n_0_26));
   NAND2_X1 i_0_0_170 (.A1(n_0_0_139), .A2(temp2[19]), .ZN(n_0_0_114));
   INV_X1 i_0_0_171 (.A(data2[19]), .ZN(n_0_0_115));
   OAI21_X1 i_0_0_172 (.A(n_0_0_116), .B1(n_0_0_117), .B2(n_0_0_139), .ZN(n_0_25));
   NAND2_X1 i_0_0_173 (.A1(n_0_0_139), .A2(temp2[20]), .ZN(n_0_0_116));
   INV_X1 i_0_0_174 (.A(data2[20]), .ZN(n_0_0_117));
   OAI21_X1 i_0_0_175 (.A(n_0_0_118), .B1(n_0_0_119), .B2(n_0_0_139), .ZN(n_0_24));
   NAND2_X1 i_0_0_176 (.A1(n_0_0_139), .A2(temp2[21]), .ZN(n_0_0_118));
   INV_X1 i_0_0_177 (.A(data2[21]), .ZN(n_0_0_119));
   OAI21_X1 i_0_0_178 (.A(n_0_0_120), .B1(n_0_0_121), .B2(n_0_0_139), .ZN(n_0_23));
   NAND2_X1 i_0_0_179 (.A1(n_0_0_139), .A2(temp2[22]), .ZN(n_0_0_120));
   INV_X1 i_0_0_180 (.A(data2[22]), .ZN(n_0_0_121));
   OAI21_X1 i_0_0_181 (.A(n_0_0_122), .B1(n_0_0_123), .B2(n_0_0_139), .ZN(n_0_22));
   NAND2_X1 i_0_0_182 (.A1(n_0_0_139), .A2(temp2[23]), .ZN(n_0_0_122));
   INV_X1 i_0_0_183 (.A(data2[23]), .ZN(n_0_0_123));
   OAI21_X1 i_0_0_184 (.A(n_0_0_124), .B1(n_0_0_125), .B2(n_0_0_139), .ZN(n_0_21));
   NAND2_X1 i_0_0_185 (.A1(n_0_0_139), .A2(temp2[24]), .ZN(n_0_0_124));
   INV_X1 i_0_0_186 (.A(data2[24]), .ZN(n_0_0_125));
   OAI21_X1 i_0_0_187 (.A(n_0_0_126), .B1(n_0_0_127), .B2(n_0_0_139), .ZN(n_0_20));
   NAND2_X1 i_0_0_188 (.A1(n_0_0_139), .A2(temp2[25]), .ZN(n_0_0_126));
   INV_X1 i_0_0_189 (.A(data2[25]), .ZN(n_0_0_127));
   OAI21_X1 i_0_0_190 (.A(n_0_0_128), .B1(n_0_0_129), .B2(n_0_0_139), .ZN(n_0_19));
   NAND2_X1 i_0_0_191 (.A1(n_0_0_139), .A2(temp2[26]), .ZN(n_0_0_128));
   INV_X1 i_0_0_192 (.A(data2[26]), .ZN(n_0_0_129));
   OAI21_X1 i_0_0_193 (.A(n_0_0_130), .B1(n_0_0_131), .B2(n_0_0_139), .ZN(n_0_18));
   NAND2_X1 i_0_0_194 (.A1(n_0_0_139), .A2(temp2[27]), .ZN(n_0_0_130));
   INV_X1 i_0_0_195 (.A(data2[27]), .ZN(n_0_0_131));
   OAI21_X1 i_0_0_196 (.A(n_0_0_132), .B1(n_0_0_133), .B2(n_0_0_139), .ZN(n_0_17));
   NAND2_X1 i_0_0_197 (.A1(n_0_0_139), .A2(temp2[28]), .ZN(n_0_0_132));
   INV_X1 i_0_0_198 (.A(data2[28]), .ZN(n_0_0_133));
   OAI21_X1 i_0_0_199 (.A(n_0_0_134), .B1(n_0_0_135), .B2(n_0_0_139), .ZN(n_0_16));
   NAND2_X1 i_0_0_200 (.A1(n_0_0_139), .A2(temp2[29]), .ZN(n_0_0_134));
   INV_X1 i_0_0_201 (.A(data2[29]), .ZN(n_0_0_135));
   OAI21_X1 i_0_0_202 (.A(n_0_0_136), .B1(n_0_0_137), .B2(n_0_0_139), .ZN(n_0_15));
   NAND2_X1 i_0_0_203 (.A1(n_0_0_139), .A2(temp2[30]), .ZN(n_0_0_136));
   INV_X1 i_0_0_204 (.A(data2[30]), .ZN(n_0_0_137));
   OAI21_X1 i_0_0_205 (.A(n_0_0_138), .B1(n_0_0_142), .B2(n_0_0_139), .ZN(n_0_14));
   NAND2_X1 i_0_0_206 (.A1(n_0_0_139), .A2(temp2[31]), .ZN(n_0_0_138));
   NAND3_X1 i_0_0_207 (.A1(n_0_8), .A2(store2), .A3(n_0_0_140), .ZN(n_0_0_139));
   NAND2_X1 i_0_0_208 (.A1(counter), .A2(n_0_0_141), .ZN(n_0_0_140));
   INV_X1 i_0_0_209 (.A(wait2), .ZN(n_0_0_141));
   INV_X1 i_0_0_210 (.A(data2[31]), .ZN(n_0_0_142));
   NAND3_X1 i_0_0_211 (.A1(n_0_0_143), .A2(n_0_0_5), .A3(n_0_0_2), .ZN(n_0_11));
   NAND3_X1 i_0_0_212 (.A1(n_0_0_6), .A2(n_0_0_3), .A3(select[0]), .ZN(n_0_0_143));
   NAND3_X1 i_0_0_213 (.A1(n_0_0_4), .A2(n_0_0_3), .A3(n_0_0_2), .ZN(n_0_12));
   NAND3_X1 i_0_0_214 (.A1(n_0_8), .A2(counter), .A3(wait2), .ZN(n_0_0_2));
   NAND3_X1 i_0_0_215 (.A1(n_0_8), .A2(n_0_13), .A3(wait1), .ZN(n_0_0_3));
   NAND3_X1 i_0_0_216 (.A1(n_0_0_6), .A2(n_0_0_5), .A3(select[1]), .ZN(n_0_0_4));
   NAND3_X1 i_0_0_217 (.A1(n_0_8), .A2(counter), .A3(store2), .ZN(n_0_0_5));
   NAND3_X1 i_0_0_218 (.A1(n_0_8), .A2(n_0_13), .A3(store1), .ZN(n_0_0_6));
   INV_X1 i_0_0_219 (.A(reset), .ZN(n_0_8));
   INV_X1 i_0_0_220 (.A(counter), .ZN(n_0_13));
   OAI21_X1 i_0_0_4 (.A(n_0_0_7), .B1(reset), .B2(n_0_0_8), .ZN(n_0_3));
   NAND2_X1 i_0_0_5 (.A1(reset), .A2(write), .ZN(n_0_0_7));
   NOR4_X1 i_0_0_6 (.A1(store1), .A2(wait2), .A3(store2), .A4(wait1), .ZN(
      n_0_0_8));
endmodule
